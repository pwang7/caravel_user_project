magic
tech sky130A
magscale 1 2
timestamp 1623917876
<< obsli1 >>
rect 1104 1377 260084 261137
<< obsm1 >>
rect 198 1368 260898 261168
<< metal2 >>
rect 1122 262535 1178 263335
rect 3330 262535 3386 263335
rect 5630 262535 5686 263335
rect 7930 262535 7986 263335
rect 10230 262535 10286 263335
rect 12530 262535 12586 263335
rect 14830 262535 14886 263335
rect 17130 262535 17186 263335
rect 19430 262535 19486 263335
rect 21730 262535 21786 263335
rect 24030 262535 24086 263335
rect 26238 262535 26294 263335
rect 28538 262535 28594 263335
rect 30838 262535 30894 263335
rect 33138 262535 33194 263335
rect 35438 262535 35494 263335
rect 37738 262535 37794 263335
rect 40038 262535 40094 263335
rect 42338 262535 42394 263335
rect 44638 262535 44694 263335
rect 46938 262535 46994 263335
rect 49146 262535 49202 263335
rect 51446 262535 51502 263335
rect 53746 262535 53802 263335
rect 56046 262535 56102 263335
rect 58346 262535 58402 263335
rect 60646 262535 60702 263335
rect 62946 262535 63002 263335
rect 65246 262535 65302 263335
rect 67546 262535 67602 263335
rect 69846 262535 69902 263335
rect 72146 262535 72202 263335
rect 74354 262535 74410 263335
rect 76654 262535 76710 263335
rect 78954 262535 79010 263335
rect 81254 262535 81310 263335
rect 83554 262535 83610 263335
rect 85854 262535 85910 263335
rect 88154 262535 88210 263335
rect 90454 262535 90510 263335
rect 92754 262535 92810 263335
rect 95054 262535 95110 263335
rect 97262 262535 97318 263335
rect 99562 262535 99618 263335
rect 101862 262535 101918 263335
rect 104162 262535 104218 263335
rect 106462 262535 106518 263335
rect 108762 262535 108818 263335
rect 111062 262535 111118 263335
rect 113362 262535 113418 263335
rect 115662 262535 115718 263335
rect 117962 262535 118018 263335
rect 120170 262535 120226 263335
rect 122470 262535 122526 263335
rect 124770 262535 124826 263335
rect 127070 262535 127126 263335
rect 129370 262535 129426 263335
rect 131670 262535 131726 263335
rect 133970 262535 134026 263335
rect 136270 262535 136326 263335
rect 138570 262535 138626 263335
rect 140870 262535 140926 263335
rect 143170 262535 143226 263335
rect 145378 262535 145434 263335
rect 147678 262535 147734 263335
rect 149978 262535 150034 263335
rect 152278 262535 152334 263335
rect 154578 262535 154634 263335
rect 156878 262535 156934 263335
rect 159178 262535 159234 263335
rect 161478 262535 161534 263335
rect 163778 262535 163834 263335
rect 166078 262535 166134 263335
rect 168286 262535 168342 263335
rect 170586 262535 170642 263335
rect 172886 262535 172942 263335
rect 175186 262535 175242 263335
rect 177486 262535 177542 263335
rect 179786 262535 179842 263335
rect 182086 262535 182142 263335
rect 184386 262535 184442 263335
rect 186686 262535 186742 263335
rect 188986 262535 189042 263335
rect 191194 262535 191250 263335
rect 193494 262535 193550 263335
rect 195794 262535 195850 263335
rect 198094 262535 198150 263335
rect 200394 262535 200450 263335
rect 202694 262535 202750 263335
rect 204994 262535 205050 263335
rect 207294 262535 207350 263335
rect 209594 262535 209650 263335
rect 211894 262535 211950 263335
rect 214194 262535 214250 263335
rect 216402 262535 216458 263335
rect 218702 262535 218758 263335
rect 221002 262535 221058 263335
rect 223302 262535 223358 263335
rect 225602 262535 225658 263335
rect 227902 262535 227958 263335
rect 230202 262535 230258 263335
rect 232502 262535 232558 263335
rect 234802 262535 234858 263335
rect 237102 262535 237158 263335
rect 239310 262535 239366 263335
rect 241610 262535 241666 263335
rect 243910 262535 243966 263335
rect 246210 262535 246266 263335
rect 248510 262535 248566 263335
rect 250810 262535 250866 263335
rect 253110 262535 253166 263335
rect 255410 262535 255466 263335
rect 257710 262535 257766 263335
rect 260010 262535 260066 263335
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3330 0 3386 800
rect 3882 0 3938 800
rect 4434 0 4490 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5998 0 6054 800
rect 6550 0 6606 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12898 0 12954 800
rect 13450 0 13506 800
rect 14002 0 14058 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21454 0 21510 800
rect 22006 0 22062 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24582 0 24638 800
rect 25134 0 25190 800
rect 25686 0 25742 800
rect 26238 0 26294 800
rect 26790 0 26846 800
rect 27250 0 27306 800
rect 27802 0 27858 800
rect 28354 0 28410 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30470 0 30526 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32034 0 32090 800
rect 32586 0 32642 800
rect 33138 0 33194 800
rect 33690 0 33746 800
rect 34242 0 34298 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39486 0 39542 800
rect 40038 0 40094 800
rect 40590 0 40646 800
rect 41142 0 41198 800
rect 41694 0 41750 800
rect 42154 0 42210 800
rect 42706 0 42762 800
rect 43258 0 43314 800
rect 43810 0 43866 800
rect 44270 0 44326 800
rect 44822 0 44878 800
rect 45374 0 45430 800
rect 45926 0 45982 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 48042 0 48098 800
rect 48594 0 48650 800
rect 49054 0 49110 800
rect 49606 0 49662 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51262 0 51318 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 53838 0 53894 800
rect 54390 0 54446 800
rect 54942 0 54998 800
rect 55494 0 55550 800
rect 56046 0 56102 800
rect 56506 0 56562 800
rect 57058 0 57114 800
rect 57610 0 57666 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59726 0 59782 800
rect 60278 0 60334 800
rect 60830 0 60886 800
rect 61290 0 61346 800
rect 61842 0 61898 800
rect 62394 0 62450 800
rect 62946 0 63002 800
rect 63498 0 63554 800
rect 63958 0 64014 800
rect 64510 0 64566 800
rect 65062 0 65118 800
rect 65614 0 65670 800
rect 66074 0 66130 800
rect 66626 0 66682 800
rect 67178 0 67234 800
rect 67730 0 67786 800
rect 68282 0 68338 800
rect 68742 0 68798 800
rect 69294 0 69350 800
rect 69846 0 69902 800
rect 70398 0 70454 800
rect 70950 0 71006 800
rect 71410 0 71466 800
rect 71962 0 72018 800
rect 72514 0 72570 800
rect 73066 0 73122 800
rect 73526 0 73582 800
rect 74078 0 74134 800
rect 74630 0 74686 800
rect 75182 0 75238 800
rect 75734 0 75790 800
rect 76194 0 76250 800
rect 76746 0 76802 800
rect 77298 0 77354 800
rect 77850 0 77906 800
rect 78310 0 78366 800
rect 78862 0 78918 800
rect 79414 0 79470 800
rect 79966 0 80022 800
rect 80518 0 80574 800
rect 80978 0 81034 800
rect 81530 0 81586 800
rect 82082 0 82138 800
rect 82634 0 82690 800
rect 83186 0 83242 800
rect 83646 0 83702 800
rect 84198 0 84254 800
rect 84750 0 84806 800
rect 85302 0 85358 800
rect 85762 0 85818 800
rect 86314 0 86370 800
rect 86866 0 86922 800
rect 87418 0 87474 800
rect 87970 0 88026 800
rect 88430 0 88486 800
rect 88982 0 89038 800
rect 89534 0 89590 800
rect 90086 0 90142 800
rect 90546 0 90602 800
rect 91098 0 91154 800
rect 91650 0 91706 800
rect 92202 0 92258 800
rect 92754 0 92810 800
rect 93214 0 93270 800
rect 93766 0 93822 800
rect 94318 0 94374 800
rect 94870 0 94926 800
rect 95330 0 95386 800
rect 95882 0 95938 800
rect 96434 0 96490 800
rect 96986 0 97042 800
rect 97538 0 97594 800
rect 97998 0 98054 800
rect 98550 0 98606 800
rect 99102 0 99158 800
rect 99654 0 99710 800
rect 100206 0 100262 800
rect 100666 0 100722 800
rect 101218 0 101274 800
rect 101770 0 101826 800
rect 102322 0 102378 800
rect 102782 0 102838 800
rect 103334 0 103390 800
rect 103886 0 103942 800
rect 104438 0 104494 800
rect 104990 0 105046 800
rect 105450 0 105506 800
rect 106002 0 106058 800
rect 106554 0 106610 800
rect 107106 0 107162 800
rect 107566 0 107622 800
rect 108118 0 108174 800
rect 108670 0 108726 800
rect 109222 0 109278 800
rect 109774 0 109830 800
rect 110234 0 110290 800
rect 110786 0 110842 800
rect 111338 0 111394 800
rect 111890 0 111946 800
rect 112442 0 112498 800
rect 112902 0 112958 800
rect 113454 0 113510 800
rect 114006 0 114062 800
rect 114558 0 114614 800
rect 115018 0 115074 800
rect 115570 0 115626 800
rect 116122 0 116178 800
rect 116674 0 116730 800
rect 117226 0 117282 800
rect 117686 0 117742 800
rect 118238 0 118294 800
rect 118790 0 118846 800
rect 119342 0 119398 800
rect 119802 0 119858 800
rect 120354 0 120410 800
rect 120906 0 120962 800
rect 121458 0 121514 800
rect 122010 0 122066 800
rect 122470 0 122526 800
rect 123022 0 123078 800
rect 123574 0 123630 800
rect 124126 0 124182 800
rect 124678 0 124734 800
rect 125138 0 125194 800
rect 125690 0 125746 800
rect 126242 0 126298 800
rect 126794 0 126850 800
rect 127254 0 127310 800
rect 127806 0 127862 800
rect 128358 0 128414 800
rect 128910 0 128966 800
rect 129462 0 129518 800
rect 129922 0 129978 800
rect 130474 0 130530 800
rect 131026 0 131082 800
rect 131578 0 131634 800
rect 132038 0 132094 800
rect 132590 0 132646 800
rect 133142 0 133198 800
rect 133694 0 133750 800
rect 134246 0 134302 800
rect 134706 0 134762 800
rect 135258 0 135314 800
rect 135810 0 135866 800
rect 136362 0 136418 800
rect 136822 0 136878 800
rect 137374 0 137430 800
rect 137926 0 137982 800
rect 138478 0 138534 800
rect 139030 0 139086 800
rect 139490 0 139546 800
rect 140042 0 140098 800
rect 140594 0 140650 800
rect 141146 0 141202 800
rect 141698 0 141754 800
rect 142158 0 142214 800
rect 142710 0 142766 800
rect 143262 0 143318 800
rect 143814 0 143870 800
rect 144274 0 144330 800
rect 144826 0 144882 800
rect 145378 0 145434 800
rect 145930 0 145986 800
rect 146482 0 146538 800
rect 146942 0 146998 800
rect 147494 0 147550 800
rect 148046 0 148102 800
rect 148598 0 148654 800
rect 149058 0 149114 800
rect 149610 0 149666 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151266 0 151322 800
rect 151726 0 151782 800
rect 152278 0 152334 800
rect 152830 0 152886 800
rect 153382 0 153438 800
rect 153934 0 153990 800
rect 154394 0 154450 800
rect 154946 0 155002 800
rect 155498 0 155554 800
rect 156050 0 156106 800
rect 156510 0 156566 800
rect 157062 0 157118 800
rect 157614 0 157670 800
rect 158166 0 158222 800
rect 158718 0 158774 800
rect 159178 0 159234 800
rect 159730 0 159786 800
rect 160282 0 160338 800
rect 160834 0 160890 800
rect 161294 0 161350 800
rect 161846 0 161902 800
rect 162398 0 162454 800
rect 162950 0 163006 800
rect 163502 0 163558 800
rect 163962 0 164018 800
rect 164514 0 164570 800
rect 165066 0 165122 800
rect 165618 0 165674 800
rect 166170 0 166226 800
rect 166630 0 166686 800
rect 167182 0 167238 800
rect 167734 0 167790 800
rect 168286 0 168342 800
rect 168746 0 168802 800
rect 169298 0 169354 800
rect 169850 0 169906 800
rect 170402 0 170458 800
rect 170954 0 171010 800
rect 171414 0 171470 800
rect 171966 0 172022 800
rect 172518 0 172574 800
rect 173070 0 173126 800
rect 173530 0 173586 800
rect 174082 0 174138 800
rect 174634 0 174690 800
rect 175186 0 175242 800
rect 175738 0 175794 800
rect 176198 0 176254 800
rect 176750 0 176806 800
rect 177302 0 177358 800
rect 177854 0 177910 800
rect 178314 0 178370 800
rect 178866 0 178922 800
rect 179418 0 179474 800
rect 179970 0 180026 800
rect 180522 0 180578 800
rect 180982 0 181038 800
rect 181534 0 181590 800
rect 182086 0 182142 800
rect 182638 0 182694 800
rect 183190 0 183246 800
rect 183650 0 183706 800
rect 184202 0 184258 800
rect 184754 0 184810 800
rect 185306 0 185362 800
rect 185766 0 185822 800
rect 186318 0 186374 800
rect 186870 0 186926 800
rect 187422 0 187478 800
rect 187974 0 188030 800
rect 188434 0 188490 800
rect 188986 0 189042 800
rect 189538 0 189594 800
rect 190090 0 190146 800
rect 190550 0 190606 800
rect 191102 0 191158 800
rect 191654 0 191710 800
rect 192206 0 192262 800
rect 192758 0 192814 800
rect 193218 0 193274 800
rect 193770 0 193826 800
rect 194322 0 194378 800
rect 194874 0 194930 800
rect 195426 0 195482 800
rect 195886 0 195942 800
rect 196438 0 196494 800
rect 196990 0 197046 800
rect 197542 0 197598 800
rect 198002 0 198058 800
rect 198554 0 198610 800
rect 199106 0 199162 800
rect 199658 0 199714 800
rect 200210 0 200266 800
rect 200670 0 200726 800
rect 201222 0 201278 800
rect 201774 0 201830 800
rect 202326 0 202382 800
rect 202786 0 202842 800
rect 203338 0 203394 800
rect 203890 0 203946 800
rect 204442 0 204498 800
rect 204994 0 205050 800
rect 205454 0 205510 800
rect 206006 0 206062 800
rect 206558 0 206614 800
rect 207110 0 207166 800
rect 207662 0 207718 800
rect 208122 0 208178 800
rect 208674 0 208730 800
rect 209226 0 209282 800
rect 209778 0 209834 800
rect 210238 0 210294 800
rect 210790 0 210846 800
rect 211342 0 211398 800
rect 211894 0 211950 800
rect 212446 0 212502 800
rect 212906 0 212962 800
rect 213458 0 213514 800
rect 214010 0 214066 800
rect 214562 0 214618 800
rect 215022 0 215078 800
rect 215574 0 215630 800
rect 216126 0 216182 800
rect 216678 0 216734 800
rect 217230 0 217286 800
rect 217690 0 217746 800
rect 218242 0 218298 800
rect 218794 0 218850 800
rect 219346 0 219402 800
rect 219806 0 219862 800
rect 220358 0 220414 800
rect 220910 0 220966 800
rect 221462 0 221518 800
rect 222014 0 222070 800
rect 222474 0 222530 800
rect 223026 0 223082 800
rect 223578 0 223634 800
rect 224130 0 224186 800
rect 224682 0 224738 800
rect 225142 0 225198 800
rect 225694 0 225750 800
rect 226246 0 226302 800
rect 226798 0 226854 800
rect 227258 0 227314 800
rect 227810 0 227866 800
rect 228362 0 228418 800
rect 228914 0 228970 800
rect 229466 0 229522 800
rect 229926 0 229982 800
rect 230478 0 230534 800
rect 231030 0 231086 800
rect 231582 0 231638 800
rect 232042 0 232098 800
rect 232594 0 232650 800
rect 233146 0 233202 800
rect 233698 0 233754 800
rect 234250 0 234306 800
rect 234710 0 234766 800
rect 235262 0 235318 800
rect 235814 0 235870 800
rect 236366 0 236422 800
rect 236918 0 236974 800
rect 237378 0 237434 800
rect 237930 0 237986 800
rect 238482 0 238538 800
rect 239034 0 239090 800
rect 239494 0 239550 800
rect 240046 0 240102 800
rect 240598 0 240654 800
rect 241150 0 241206 800
rect 241702 0 241758 800
rect 242162 0 242218 800
rect 242714 0 242770 800
rect 243266 0 243322 800
rect 243818 0 243874 800
rect 244278 0 244334 800
rect 244830 0 244886 800
rect 245382 0 245438 800
rect 245934 0 245990 800
rect 246486 0 246542 800
rect 246946 0 247002 800
rect 247498 0 247554 800
rect 248050 0 248106 800
rect 248602 0 248658 800
rect 249154 0 249210 800
rect 249614 0 249670 800
rect 250166 0 250222 800
rect 250718 0 250774 800
rect 251270 0 251326 800
rect 251730 0 251786 800
rect 252282 0 252338 800
rect 252834 0 252890 800
rect 253386 0 253442 800
rect 253938 0 253994 800
rect 254398 0 254454 800
rect 254950 0 255006 800
rect 255502 0 255558 800
rect 256054 0 256110 800
rect 256514 0 256570 800
rect 257066 0 257122 800
rect 257618 0 257674 800
rect 258170 0 258226 800
rect 258722 0 258778 800
rect 259182 0 259238 800
rect 259734 0 259790 800
rect 260286 0 260342 800
rect 260838 0 260894 800
<< obsm2 >>
rect 204 262479 1066 262535
rect 1234 262479 3274 262535
rect 3442 262479 5574 262535
rect 5742 262479 7874 262535
rect 8042 262479 10174 262535
rect 10342 262479 12474 262535
rect 12642 262479 14774 262535
rect 14942 262479 17074 262535
rect 17242 262479 19374 262535
rect 19542 262479 21674 262535
rect 21842 262479 23974 262535
rect 24142 262479 26182 262535
rect 26350 262479 28482 262535
rect 28650 262479 30782 262535
rect 30950 262479 33082 262535
rect 33250 262479 35382 262535
rect 35550 262479 37682 262535
rect 37850 262479 39982 262535
rect 40150 262479 42282 262535
rect 42450 262479 44582 262535
rect 44750 262479 46882 262535
rect 47050 262479 49090 262535
rect 49258 262479 51390 262535
rect 51558 262479 53690 262535
rect 53858 262479 55990 262535
rect 56158 262479 58290 262535
rect 58458 262479 60590 262535
rect 60758 262479 62890 262535
rect 63058 262479 65190 262535
rect 65358 262479 67490 262535
rect 67658 262479 69790 262535
rect 69958 262479 72090 262535
rect 72258 262479 74298 262535
rect 74466 262479 76598 262535
rect 76766 262479 78898 262535
rect 79066 262479 81198 262535
rect 81366 262479 83498 262535
rect 83666 262479 85798 262535
rect 85966 262479 88098 262535
rect 88266 262479 90398 262535
rect 90566 262479 92698 262535
rect 92866 262479 94998 262535
rect 95166 262479 97206 262535
rect 97374 262479 99506 262535
rect 99674 262479 101806 262535
rect 101974 262479 104106 262535
rect 104274 262479 106406 262535
rect 106574 262479 108706 262535
rect 108874 262479 111006 262535
rect 111174 262479 113306 262535
rect 113474 262479 115606 262535
rect 115774 262479 117906 262535
rect 118074 262479 120114 262535
rect 120282 262479 122414 262535
rect 122582 262479 124714 262535
rect 124882 262479 127014 262535
rect 127182 262479 129314 262535
rect 129482 262479 131614 262535
rect 131782 262479 133914 262535
rect 134082 262479 136214 262535
rect 136382 262479 138514 262535
rect 138682 262479 140814 262535
rect 140982 262479 143114 262535
rect 143282 262479 145322 262535
rect 145490 262479 147622 262535
rect 147790 262479 149922 262535
rect 150090 262479 152222 262535
rect 152390 262479 154522 262535
rect 154690 262479 156822 262535
rect 156990 262479 159122 262535
rect 159290 262479 161422 262535
rect 161590 262479 163722 262535
rect 163890 262479 166022 262535
rect 166190 262479 168230 262535
rect 168398 262479 170530 262535
rect 170698 262479 172830 262535
rect 172998 262479 175130 262535
rect 175298 262479 177430 262535
rect 177598 262479 179730 262535
rect 179898 262479 182030 262535
rect 182198 262479 184330 262535
rect 184498 262479 186630 262535
rect 186798 262479 188930 262535
rect 189098 262479 191138 262535
rect 191306 262479 193438 262535
rect 193606 262479 195738 262535
rect 195906 262479 198038 262535
rect 198206 262479 200338 262535
rect 200506 262479 202638 262535
rect 202806 262479 204938 262535
rect 205106 262479 207238 262535
rect 207406 262479 209538 262535
rect 209706 262479 211838 262535
rect 212006 262479 214138 262535
rect 214306 262479 216346 262535
rect 216514 262479 218646 262535
rect 218814 262479 220946 262535
rect 221114 262479 223246 262535
rect 223414 262479 225546 262535
rect 225714 262479 227846 262535
rect 228014 262479 230146 262535
rect 230314 262479 232446 262535
rect 232614 262479 234746 262535
rect 234914 262479 237046 262535
rect 237214 262479 239254 262535
rect 239422 262479 241554 262535
rect 241722 262479 243854 262535
rect 244022 262479 246154 262535
rect 246322 262479 248454 262535
rect 248622 262479 250754 262535
rect 250922 262479 253054 262535
rect 253222 262479 255354 262535
rect 255522 262479 257654 262535
rect 257822 262479 259954 262535
rect 260122 262479 260892 262535
rect 204 856 260892 262479
rect 314 800 606 856
rect 774 800 1158 856
rect 1326 800 1710 856
rect 1878 800 2262 856
rect 2430 800 2722 856
rect 2890 800 3274 856
rect 3442 800 3826 856
rect 3994 800 4378 856
rect 4546 800 4930 856
rect 5098 800 5390 856
rect 5558 800 5942 856
rect 6110 800 6494 856
rect 6662 800 7046 856
rect 7214 800 7506 856
rect 7674 800 8058 856
rect 8226 800 8610 856
rect 8778 800 9162 856
rect 9330 800 9714 856
rect 9882 800 10174 856
rect 10342 800 10726 856
rect 10894 800 11278 856
rect 11446 800 11830 856
rect 11998 800 12290 856
rect 12458 800 12842 856
rect 13010 800 13394 856
rect 13562 800 13946 856
rect 14114 800 14498 856
rect 14666 800 14958 856
rect 15126 800 15510 856
rect 15678 800 16062 856
rect 16230 800 16614 856
rect 16782 800 17166 856
rect 17334 800 17626 856
rect 17794 800 18178 856
rect 18346 800 18730 856
rect 18898 800 19282 856
rect 19450 800 19742 856
rect 19910 800 20294 856
rect 20462 800 20846 856
rect 21014 800 21398 856
rect 21566 800 21950 856
rect 22118 800 22410 856
rect 22578 800 22962 856
rect 23130 800 23514 856
rect 23682 800 24066 856
rect 24234 800 24526 856
rect 24694 800 25078 856
rect 25246 800 25630 856
rect 25798 800 26182 856
rect 26350 800 26734 856
rect 26902 800 27194 856
rect 27362 800 27746 856
rect 27914 800 28298 856
rect 28466 800 28850 856
rect 29018 800 29402 856
rect 29570 800 29862 856
rect 30030 800 30414 856
rect 30582 800 30966 856
rect 31134 800 31518 856
rect 31686 800 31978 856
rect 32146 800 32530 856
rect 32698 800 33082 856
rect 33250 800 33634 856
rect 33802 800 34186 856
rect 34354 800 34646 856
rect 34814 800 35198 856
rect 35366 800 35750 856
rect 35918 800 36302 856
rect 36470 800 36762 856
rect 36930 800 37314 856
rect 37482 800 37866 856
rect 38034 800 38418 856
rect 38586 800 38970 856
rect 39138 800 39430 856
rect 39598 800 39982 856
rect 40150 800 40534 856
rect 40702 800 41086 856
rect 41254 800 41638 856
rect 41806 800 42098 856
rect 42266 800 42650 856
rect 42818 800 43202 856
rect 43370 800 43754 856
rect 43922 800 44214 856
rect 44382 800 44766 856
rect 44934 800 45318 856
rect 45486 800 45870 856
rect 46038 800 46422 856
rect 46590 800 46882 856
rect 47050 800 47434 856
rect 47602 800 47986 856
rect 48154 800 48538 856
rect 48706 800 48998 856
rect 49166 800 49550 856
rect 49718 800 50102 856
rect 50270 800 50654 856
rect 50822 800 51206 856
rect 51374 800 51666 856
rect 51834 800 52218 856
rect 52386 800 52770 856
rect 52938 800 53322 856
rect 53490 800 53782 856
rect 53950 800 54334 856
rect 54502 800 54886 856
rect 55054 800 55438 856
rect 55606 800 55990 856
rect 56158 800 56450 856
rect 56618 800 57002 856
rect 57170 800 57554 856
rect 57722 800 58106 856
rect 58274 800 58658 856
rect 58826 800 59118 856
rect 59286 800 59670 856
rect 59838 800 60222 856
rect 60390 800 60774 856
rect 60942 800 61234 856
rect 61402 800 61786 856
rect 61954 800 62338 856
rect 62506 800 62890 856
rect 63058 800 63442 856
rect 63610 800 63902 856
rect 64070 800 64454 856
rect 64622 800 65006 856
rect 65174 800 65558 856
rect 65726 800 66018 856
rect 66186 800 66570 856
rect 66738 800 67122 856
rect 67290 800 67674 856
rect 67842 800 68226 856
rect 68394 800 68686 856
rect 68854 800 69238 856
rect 69406 800 69790 856
rect 69958 800 70342 856
rect 70510 800 70894 856
rect 71062 800 71354 856
rect 71522 800 71906 856
rect 72074 800 72458 856
rect 72626 800 73010 856
rect 73178 800 73470 856
rect 73638 800 74022 856
rect 74190 800 74574 856
rect 74742 800 75126 856
rect 75294 800 75678 856
rect 75846 800 76138 856
rect 76306 800 76690 856
rect 76858 800 77242 856
rect 77410 800 77794 856
rect 77962 800 78254 856
rect 78422 800 78806 856
rect 78974 800 79358 856
rect 79526 800 79910 856
rect 80078 800 80462 856
rect 80630 800 80922 856
rect 81090 800 81474 856
rect 81642 800 82026 856
rect 82194 800 82578 856
rect 82746 800 83130 856
rect 83298 800 83590 856
rect 83758 800 84142 856
rect 84310 800 84694 856
rect 84862 800 85246 856
rect 85414 800 85706 856
rect 85874 800 86258 856
rect 86426 800 86810 856
rect 86978 800 87362 856
rect 87530 800 87914 856
rect 88082 800 88374 856
rect 88542 800 88926 856
rect 89094 800 89478 856
rect 89646 800 90030 856
rect 90198 800 90490 856
rect 90658 800 91042 856
rect 91210 800 91594 856
rect 91762 800 92146 856
rect 92314 800 92698 856
rect 92866 800 93158 856
rect 93326 800 93710 856
rect 93878 800 94262 856
rect 94430 800 94814 856
rect 94982 800 95274 856
rect 95442 800 95826 856
rect 95994 800 96378 856
rect 96546 800 96930 856
rect 97098 800 97482 856
rect 97650 800 97942 856
rect 98110 800 98494 856
rect 98662 800 99046 856
rect 99214 800 99598 856
rect 99766 800 100150 856
rect 100318 800 100610 856
rect 100778 800 101162 856
rect 101330 800 101714 856
rect 101882 800 102266 856
rect 102434 800 102726 856
rect 102894 800 103278 856
rect 103446 800 103830 856
rect 103998 800 104382 856
rect 104550 800 104934 856
rect 105102 800 105394 856
rect 105562 800 105946 856
rect 106114 800 106498 856
rect 106666 800 107050 856
rect 107218 800 107510 856
rect 107678 800 108062 856
rect 108230 800 108614 856
rect 108782 800 109166 856
rect 109334 800 109718 856
rect 109886 800 110178 856
rect 110346 800 110730 856
rect 110898 800 111282 856
rect 111450 800 111834 856
rect 112002 800 112386 856
rect 112554 800 112846 856
rect 113014 800 113398 856
rect 113566 800 113950 856
rect 114118 800 114502 856
rect 114670 800 114962 856
rect 115130 800 115514 856
rect 115682 800 116066 856
rect 116234 800 116618 856
rect 116786 800 117170 856
rect 117338 800 117630 856
rect 117798 800 118182 856
rect 118350 800 118734 856
rect 118902 800 119286 856
rect 119454 800 119746 856
rect 119914 800 120298 856
rect 120466 800 120850 856
rect 121018 800 121402 856
rect 121570 800 121954 856
rect 122122 800 122414 856
rect 122582 800 122966 856
rect 123134 800 123518 856
rect 123686 800 124070 856
rect 124238 800 124622 856
rect 124790 800 125082 856
rect 125250 800 125634 856
rect 125802 800 126186 856
rect 126354 800 126738 856
rect 126906 800 127198 856
rect 127366 800 127750 856
rect 127918 800 128302 856
rect 128470 800 128854 856
rect 129022 800 129406 856
rect 129574 800 129866 856
rect 130034 800 130418 856
rect 130586 800 130970 856
rect 131138 800 131522 856
rect 131690 800 131982 856
rect 132150 800 132534 856
rect 132702 800 133086 856
rect 133254 800 133638 856
rect 133806 800 134190 856
rect 134358 800 134650 856
rect 134818 800 135202 856
rect 135370 800 135754 856
rect 135922 800 136306 856
rect 136474 800 136766 856
rect 136934 800 137318 856
rect 137486 800 137870 856
rect 138038 800 138422 856
rect 138590 800 138974 856
rect 139142 800 139434 856
rect 139602 800 139986 856
rect 140154 800 140538 856
rect 140706 800 141090 856
rect 141258 800 141642 856
rect 141810 800 142102 856
rect 142270 800 142654 856
rect 142822 800 143206 856
rect 143374 800 143758 856
rect 143926 800 144218 856
rect 144386 800 144770 856
rect 144938 800 145322 856
rect 145490 800 145874 856
rect 146042 800 146426 856
rect 146594 800 146886 856
rect 147054 800 147438 856
rect 147606 800 147990 856
rect 148158 800 148542 856
rect 148710 800 149002 856
rect 149170 800 149554 856
rect 149722 800 150106 856
rect 150274 800 150658 856
rect 150826 800 151210 856
rect 151378 800 151670 856
rect 151838 800 152222 856
rect 152390 800 152774 856
rect 152942 800 153326 856
rect 153494 800 153878 856
rect 154046 800 154338 856
rect 154506 800 154890 856
rect 155058 800 155442 856
rect 155610 800 155994 856
rect 156162 800 156454 856
rect 156622 800 157006 856
rect 157174 800 157558 856
rect 157726 800 158110 856
rect 158278 800 158662 856
rect 158830 800 159122 856
rect 159290 800 159674 856
rect 159842 800 160226 856
rect 160394 800 160778 856
rect 160946 800 161238 856
rect 161406 800 161790 856
rect 161958 800 162342 856
rect 162510 800 162894 856
rect 163062 800 163446 856
rect 163614 800 163906 856
rect 164074 800 164458 856
rect 164626 800 165010 856
rect 165178 800 165562 856
rect 165730 800 166114 856
rect 166282 800 166574 856
rect 166742 800 167126 856
rect 167294 800 167678 856
rect 167846 800 168230 856
rect 168398 800 168690 856
rect 168858 800 169242 856
rect 169410 800 169794 856
rect 169962 800 170346 856
rect 170514 800 170898 856
rect 171066 800 171358 856
rect 171526 800 171910 856
rect 172078 800 172462 856
rect 172630 800 173014 856
rect 173182 800 173474 856
rect 173642 800 174026 856
rect 174194 800 174578 856
rect 174746 800 175130 856
rect 175298 800 175682 856
rect 175850 800 176142 856
rect 176310 800 176694 856
rect 176862 800 177246 856
rect 177414 800 177798 856
rect 177966 800 178258 856
rect 178426 800 178810 856
rect 178978 800 179362 856
rect 179530 800 179914 856
rect 180082 800 180466 856
rect 180634 800 180926 856
rect 181094 800 181478 856
rect 181646 800 182030 856
rect 182198 800 182582 856
rect 182750 800 183134 856
rect 183302 800 183594 856
rect 183762 800 184146 856
rect 184314 800 184698 856
rect 184866 800 185250 856
rect 185418 800 185710 856
rect 185878 800 186262 856
rect 186430 800 186814 856
rect 186982 800 187366 856
rect 187534 800 187918 856
rect 188086 800 188378 856
rect 188546 800 188930 856
rect 189098 800 189482 856
rect 189650 800 190034 856
rect 190202 800 190494 856
rect 190662 800 191046 856
rect 191214 800 191598 856
rect 191766 800 192150 856
rect 192318 800 192702 856
rect 192870 800 193162 856
rect 193330 800 193714 856
rect 193882 800 194266 856
rect 194434 800 194818 856
rect 194986 800 195370 856
rect 195538 800 195830 856
rect 195998 800 196382 856
rect 196550 800 196934 856
rect 197102 800 197486 856
rect 197654 800 197946 856
rect 198114 800 198498 856
rect 198666 800 199050 856
rect 199218 800 199602 856
rect 199770 800 200154 856
rect 200322 800 200614 856
rect 200782 800 201166 856
rect 201334 800 201718 856
rect 201886 800 202270 856
rect 202438 800 202730 856
rect 202898 800 203282 856
rect 203450 800 203834 856
rect 204002 800 204386 856
rect 204554 800 204938 856
rect 205106 800 205398 856
rect 205566 800 205950 856
rect 206118 800 206502 856
rect 206670 800 207054 856
rect 207222 800 207606 856
rect 207774 800 208066 856
rect 208234 800 208618 856
rect 208786 800 209170 856
rect 209338 800 209722 856
rect 209890 800 210182 856
rect 210350 800 210734 856
rect 210902 800 211286 856
rect 211454 800 211838 856
rect 212006 800 212390 856
rect 212558 800 212850 856
rect 213018 800 213402 856
rect 213570 800 213954 856
rect 214122 800 214506 856
rect 214674 800 214966 856
rect 215134 800 215518 856
rect 215686 800 216070 856
rect 216238 800 216622 856
rect 216790 800 217174 856
rect 217342 800 217634 856
rect 217802 800 218186 856
rect 218354 800 218738 856
rect 218906 800 219290 856
rect 219458 800 219750 856
rect 219918 800 220302 856
rect 220470 800 220854 856
rect 221022 800 221406 856
rect 221574 800 221958 856
rect 222126 800 222418 856
rect 222586 800 222970 856
rect 223138 800 223522 856
rect 223690 800 224074 856
rect 224242 800 224626 856
rect 224794 800 225086 856
rect 225254 800 225638 856
rect 225806 800 226190 856
rect 226358 800 226742 856
rect 226910 800 227202 856
rect 227370 800 227754 856
rect 227922 800 228306 856
rect 228474 800 228858 856
rect 229026 800 229410 856
rect 229578 800 229870 856
rect 230038 800 230422 856
rect 230590 800 230974 856
rect 231142 800 231526 856
rect 231694 800 231986 856
rect 232154 800 232538 856
rect 232706 800 233090 856
rect 233258 800 233642 856
rect 233810 800 234194 856
rect 234362 800 234654 856
rect 234822 800 235206 856
rect 235374 800 235758 856
rect 235926 800 236310 856
rect 236478 800 236862 856
rect 237030 800 237322 856
rect 237490 800 237874 856
rect 238042 800 238426 856
rect 238594 800 238978 856
rect 239146 800 239438 856
rect 239606 800 239990 856
rect 240158 800 240542 856
rect 240710 800 241094 856
rect 241262 800 241646 856
rect 241814 800 242106 856
rect 242274 800 242658 856
rect 242826 800 243210 856
rect 243378 800 243762 856
rect 243930 800 244222 856
rect 244390 800 244774 856
rect 244942 800 245326 856
rect 245494 800 245878 856
rect 246046 800 246430 856
rect 246598 800 246890 856
rect 247058 800 247442 856
rect 247610 800 247994 856
rect 248162 800 248546 856
rect 248714 800 249098 856
rect 249266 800 249558 856
rect 249726 800 250110 856
rect 250278 800 250662 856
rect 250830 800 251214 856
rect 251382 800 251674 856
rect 251842 800 252226 856
rect 252394 800 252778 856
rect 252946 800 253330 856
rect 253498 800 253882 856
rect 254050 800 254342 856
rect 254510 800 254894 856
rect 255062 800 255446 856
rect 255614 800 255998 856
rect 256166 800 256458 856
rect 256626 800 257010 856
rect 257178 800 257562 856
rect 257730 800 258114 856
rect 258282 800 258666 856
rect 258834 800 259126 856
rect 259294 800 259678 856
rect 259846 800 260230 856
rect 260398 800 260782 856
<< metal3 >>
rect 0 131656 800 131776
rect 260391 131656 261191 131776
<< obsm3 >>
rect 800 131856 260391 261153
rect 880 131576 260311 131856
rect 800 2143 260391 131576
<< metal4 >>
rect 4208 2128 4528 261168
rect 4868 2176 5188 261120
rect 5528 2176 5848 261120
rect 6188 2176 6508 261120
rect 19568 2128 19888 261168
rect 20228 2176 20548 261120
rect 20888 2176 21208 261120
rect 21548 2176 21868 261120
rect 34928 2128 35248 261168
rect 35588 2176 35908 261120
rect 36248 2176 36568 261120
rect 36908 2176 37228 261120
rect 50288 2128 50608 261168
rect 50948 2176 51268 261120
rect 51608 2176 51928 261120
rect 52268 2176 52588 261120
rect 65648 2128 65968 261168
rect 66308 2176 66628 261120
rect 66968 2176 67288 261120
rect 67628 2176 67948 261120
rect 81008 2128 81328 261168
rect 81668 2176 81988 261120
rect 82328 2176 82648 261120
rect 82988 2176 83308 261120
rect 96368 2128 96688 261168
rect 97028 2176 97348 261120
rect 97688 2176 98008 261120
rect 98348 2176 98668 261120
rect 111728 2128 112048 261168
rect 112388 2176 112708 261120
rect 113048 2176 113368 261120
rect 113708 2176 114028 261120
rect 127088 2128 127408 261168
rect 127748 2176 128068 261120
rect 128408 2176 128728 261120
rect 129068 2176 129388 261120
rect 142448 2128 142768 261168
rect 143108 2176 143428 261120
rect 143768 2176 144088 261120
rect 144428 2176 144748 261120
rect 157808 2128 158128 261168
rect 158468 2176 158788 261120
rect 159128 2176 159448 261120
rect 159788 2176 160108 261120
rect 173168 2128 173488 261168
rect 173828 2176 174148 261120
rect 174488 2176 174808 261120
rect 175148 2176 175468 261120
rect 188528 2128 188848 261168
rect 189188 2176 189508 261120
rect 189848 2176 190168 261120
rect 190508 2176 190828 261120
rect 203888 2128 204208 261168
rect 204548 2176 204868 261120
rect 205208 2176 205528 261120
rect 205868 2176 206188 261120
rect 219248 2128 219568 261168
rect 219908 2176 220228 261120
rect 220568 2176 220888 261120
rect 221228 2176 221548 261120
rect 234608 2128 234928 261168
rect 235268 2176 235588 261120
rect 235928 2176 236248 261120
rect 236588 2176 236908 261120
rect 249968 2128 250288 261168
rect 250628 2176 250948 261120
rect 251288 2176 251608 261120
rect 251948 2176 252268 261120
<< obsm4 >>
rect 49923 56339 50208 212397
rect 50688 56339 50868 212397
rect 51348 56339 51528 212397
rect 52008 56339 52188 212397
rect 52668 56339 65568 212397
rect 66048 56339 66228 212397
rect 66708 56339 66888 212397
rect 67368 56339 67548 212397
rect 68028 56339 80928 212397
rect 81408 56339 81588 212397
rect 82068 56339 82248 212397
rect 82728 56339 82908 212397
rect 83388 56339 96288 212397
rect 96768 56339 96948 212397
rect 97428 56339 97608 212397
rect 98088 56339 98268 212397
rect 98748 56339 111648 212397
rect 112128 56339 112308 212397
rect 112788 56339 112968 212397
rect 113448 56339 113628 212397
rect 114108 56339 127008 212397
rect 127488 56339 127668 212397
rect 128148 56339 128328 212397
rect 128808 56339 128988 212397
rect 129468 56339 142368 212397
rect 142848 56339 143028 212397
rect 143508 56339 143688 212397
rect 144168 56339 144348 212397
rect 144828 56339 157728 212397
rect 158208 56339 158388 212397
rect 158868 56339 159048 212397
rect 159528 56339 159708 212397
rect 160188 56339 173088 212397
rect 173568 56339 173748 212397
rect 174228 56339 174408 212397
rect 174888 56339 175068 212397
rect 175548 56339 188448 212397
rect 188928 56339 189108 212397
rect 189588 56339 189768 212397
rect 190248 56339 190428 212397
rect 190908 56339 203808 212397
<< labels >>
rlabel metal2 s 1122 262535 1178 263335 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 69846 262535 69902 263335 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 76654 262535 76710 263335 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 83554 262535 83610 263335 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 90454 262535 90510 263335 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 97262 262535 97318 263335 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 104162 262535 104218 263335 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 111062 262535 111118 263335 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 117962 262535 118018 263335 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 124770 262535 124826 263335 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 131670 262535 131726 263335 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7930 262535 7986 263335 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 138570 262535 138626 263335 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 145378 262535 145434 263335 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 152278 262535 152334 263335 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 159178 262535 159234 263335 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 166078 262535 166134 263335 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 172886 262535 172942 263335 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 179786 262535 179842 263335 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 186686 262535 186742 263335 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 193494 262535 193550 263335 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 200394 262535 200450 263335 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14830 262535 14886 263335 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 207294 262535 207350 263335 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 214194 262535 214250 263335 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 221002 262535 221058 263335 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 227902 262535 227958 263335 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 234802 262535 234858 263335 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 241610 262535 241666 263335 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 248510 262535 248566 263335 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 255410 262535 255466 263335 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 21730 262535 21786 263335 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 28538 262535 28594 263335 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 35438 262535 35494 263335 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 42338 262535 42394 263335 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 49146 262535 49202 263335 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 56046 262535 56102 263335 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 62946 262535 63002 263335 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3330 262535 3386 263335 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 72146 262535 72202 263335 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 78954 262535 79010 263335 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 85854 262535 85910 263335 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 92754 262535 92810 263335 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 99562 262535 99618 263335 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 106462 262535 106518 263335 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 113362 262535 113418 263335 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 120170 262535 120226 263335 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 127070 262535 127126 263335 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 133970 262535 134026 263335 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 10230 262535 10286 263335 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 140870 262535 140926 263335 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 147678 262535 147734 263335 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 154578 262535 154634 263335 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 161478 262535 161534 263335 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 168286 262535 168342 263335 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 175186 262535 175242 263335 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 182086 262535 182142 263335 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 188986 262535 189042 263335 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 195794 262535 195850 263335 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 202694 262535 202750 263335 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 17130 262535 17186 263335 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 209594 262535 209650 263335 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 216402 262535 216458 263335 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 223302 262535 223358 263335 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 230202 262535 230258 263335 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 237102 262535 237158 263335 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 243910 262535 243966 263335 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 250810 262535 250866 263335 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 257710 262535 257766 263335 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 24030 262535 24086 263335 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 30838 262535 30894 263335 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 37738 262535 37794 263335 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 44638 262535 44694 263335 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 51446 262535 51502 263335 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 58346 262535 58402 263335 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 65246 262535 65302 263335 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5630 262535 5686 263335 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 74354 262535 74410 263335 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 81254 262535 81310 263335 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 88154 262535 88210 263335 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 95054 262535 95110 263335 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 101862 262535 101918 263335 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 108762 262535 108818 263335 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 115662 262535 115718 263335 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 122470 262535 122526 263335 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 129370 262535 129426 263335 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 136270 262535 136326 263335 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 12530 262535 12586 263335 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 143170 262535 143226 263335 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 149978 262535 150034 263335 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 156878 262535 156934 263335 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 163778 262535 163834 263335 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 170586 262535 170642 263335 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 177486 262535 177542 263335 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 184386 262535 184442 263335 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 191194 262535 191250 263335 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 198094 262535 198150 263335 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 204994 262535 205050 263335 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 19430 262535 19486 263335 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 211894 262535 211950 263335 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 218702 262535 218758 263335 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 225602 262535 225658 263335 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 232502 262535 232558 263335 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 239310 262535 239366 263335 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 246210 262535 246266 263335 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 253110 262535 253166 263335 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 260010 262535 260066 263335 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 26238 262535 26294 263335 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 33138 262535 33194 263335 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 40038 262535 40094 263335 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 46938 262535 46994 263335 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 53746 262535 53802 263335 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 60646 262535 60702 263335 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 67546 262535 67602 263335 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 260838 0 260894 800 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 260391 131656 261191 131776 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 216126 0 216182 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 217690 0 217746 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 219346 0 219402 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 232042 0 232098 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 233698 0 233754 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 238482 0 238538 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 240046 0 240102 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 243266 0 243322 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 246486 0 246542 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 248050 0 248106 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 251270 0 251326 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 252834 0 252890 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 256054 0 256110 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 163502 0 163558 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 196990 0 197046 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 200210 0 200266 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 201774 0 201830 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 211342 0 211398 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 214562 0 214618 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 216678 0 216734 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 218242 0 218298 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 219806 0 219862 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 221462 0 221518 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 223026 0 223082 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 224682 0 224738 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 226246 0 226302 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 227810 0 227866 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 229466 0 229522 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 231030 0 231086 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 232594 0 232650 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 237378 0 237434 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 239034 0 239090 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 240598 0 240654 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 242162 0 242218 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 243818 0 243874 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 246946 0 247002 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 248602 0 248658 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 250166 0 250222 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 251730 0 251786 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 253386 0 253442 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 254950 0 255006 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 256514 0 256570 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 258170 0 258226 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 259734 0 259790 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 148046 0 148102 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 151266 0 151322 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 160834 0 160890 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 162398 0 162454 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 167182 0 167238 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 170402 0 170458 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 171966 0 172022 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 179970 0 180026 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 181534 0 181590 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 184754 0 184810 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 187974 0 188030 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 189538 0 189594 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 191102 0 191158 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 192758 0 192814 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 194322 0 194378 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 195886 0 195942 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 197542 0 197598 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 200670 0 200726 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 202326 0 202382 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 203890 0 203946 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 205454 0 205510 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 207110 0 207166 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 208674 0 208730 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 210238 0 210294 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 211894 0 211950 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 213458 0 213514 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 215022 0 215078 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 217230 0 217286 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 222014 0 222070 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 234710 0 234766 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 237930 0 237986 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 239494 0 239550 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 241150 0 241206 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 242714 0 242770 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 244278 0 244334 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 245934 0 245990 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 247498 0 247554 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 249154 0 249210 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 250718 0 250774 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 252282 0 252338 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 255502 0 255558 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 257066 0 257122 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 258722 0 258778 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 260286 0 260342 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 183650 0 183706 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 191654 0 191710 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 194874 0 194930 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 204442 0 204498 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 206006 0 206062 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 209226 0 209282 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 215574 0 215630 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 249968 2128 250288 261168 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 261168 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 261168 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 261168 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 261168 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 261168 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 261168 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 261168 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 261168 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 234608 2128 234928 261168 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 261168 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 261168 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 261168 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 261168 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 261168 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 261168 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 261168 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 250628 2176 250948 261120 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 261120 6 vccd2
port 626 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 261120 6 vccd2
port 627 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 261120 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 261120 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 261120 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 261120 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 261120 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 261120 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 235268 2176 235588 261120 6 vssd2
port 634 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 261120 6 vssd2
port 635 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 261120 6 vssd2
port 636 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 261120 6 vssd2
port 637 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 261120 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 261120 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 261120 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 261120 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 251288 2176 251608 261120 6 vdda1
port 642 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 261120 6 vdda1
port 643 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 261120 6 vdda1
port 644 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 261120 6 vdda1
port 645 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 261120 6 vdda1
port 646 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 261120 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 261120 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 261120 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 261120 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 235928 2176 236248 261120 6 vssa1
port 651 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 261120 6 vssa1
port 652 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 261120 6 vssa1
port 653 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 261120 6 vssa1
port 654 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 261120 6 vssa1
port 655 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 261120 6 vssa1
port 656 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 261120 6 vssa1
port 657 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 261120 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 251948 2176 252268 261120 6 vdda2
port 659 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 261120 6 vdda2
port 660 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 261120 6 vdda2
port 661 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 261120 6 vdda2
port 662 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 261120 6 vdda2
port 663 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 261120 6 vdda2
port 664 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 261120 6 vdda2
port 665 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 261120 6 vdda2
port 666 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 261120 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 236588 2176 236908 261120 6 vssa2
port 668 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 261120 6 vssa2
port 669 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 261120 6 vssa2
port 670 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 261120 6 vssa2
port 671 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 261120 6 vssa2
port 672 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 261120 6 vssa2
port 673 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 261120 6 vssa2
port 674 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 261120 6 vssa2
port 675 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 261191 263335
string LEFview TRUE
string GDS_FILE /project/openlane/axi_dma/runs/axi_dma/results/magic/axi_dma.gds
string GDS_END 95116034
string GDS_START 1118362
<< end >>

