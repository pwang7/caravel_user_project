magic
tech sky130A
magscale 1 2
timestamp 1623396513
<< obsli1 >>
rect 1104 1309 261372 262225
<< obsm1 >>
rect 198 1300 262186 262256
<< metal2 >>
rect 1122 263849 1178 264649
rect 3330 263849 3386 264649
rect 5630 263849 5686 264649
rect 7838 263849 7894 264649
rect 10138 263849 10194 264649
rect 12346 263849 12402 264649
rect 14646 263849 14702 264649
rect 16946 263849 17002 264649
rect 19154 263849 19210 264649
rect 21454 263849 21510 264649
rect 23662 263849 23718 264649
rect 25962 263849 26018 264649
rect 28262 263849 28318 264649
rect 30470 263849 30526 264649
rect 32770 263849 32826 264649
rect 34978 263849 35034 264649
rect 37278 263849 37334 264649
rect 39578 263849 39634 264649
rect 41786 263849 41842 264649
rect 44086 263849 44142 264649
rect 46294 263849 46350 264649
rect 48594 263849 48650 264649
rect 50894 263849 50950 264649
rect 53102 263849 53158 264649
rect 55402 263849 55458 264649
rect 57610 263849 57666 264649
rect 59910 263849 59966 264649
rect 62210 263849 62266 264649
rect 64418 263849 64474 264649
rect 66718 263849 66774 264649
rect 68926 263849 68982 264649
rect 71226 263849 71282 264649
rect 73526 263849 73582 264649
rect 75734 263849 75790 264649
rect 78034 263849 78090 264649
rect 80242 263849 80298 264649
rect 82542 263849 82598 264649
rect 84842 263849 84898 264649
rect 87050 263849 87106 264649
rect 89350 263849 89406 264649
rect 91558 263849 91614 264649
rect 93858 263849 93914 264649
rect 96066 263849 96122 264649
rect 98366 263849 98422 264649
rect 100666 263849 100722 264649
rect 102874 263849 102930 264649
rect 105174 263849 105230 264649
rect 107382 263849 107438 264649
rect 109682 263849 109738 264649
rect 111982 263849 112038 264649
rect 114190 263849 114246 264649
rect 116490 263849 116546 264649
rect 118698 263849 118754 264649
rect 120998 263849 121054 264649
rect 123298 263849 123354 264649
rect 125506 263849 125562 264649
rect 127806 263849 127862 264649
rect 130014 263849 130070 264649
rect 132314 263849 132370 264649
rect 134614 263849 134670 264649
rect 136822 263849 136878 264649
rect 139122 263849 139178 264649
rect 141330 263849 141386 264649
rect 143630 263849 143686 264649
rect 145930 263849 145986 264649
rect 148138 263849 148194 264649
rect 150438 263849 150494 264649
rect 152646 263849 152702 264649
rect 154946 263849 155002 264649
rect 157246 263849 157302 264649
rect 159454 263849 159510 264649
rect 161754 263849 161810 264649
rect 163962 263849 164018 264649
rect 166262 263849 166318 264649
rect 168562 263849 168618 264649
rect 170770 263849 170826 264649
rect 173070 263849 173126 264649
rect 175278 263849 175334 264649
rect 177578 263849 177634 264649
rect 179786 263849 179842 264649
rect 182086 263849 182142 264649
rect 184386 263849 184442 264649
rect 186594 263849 186650 264649
rect 188894 263849 188950 264649
rect 191102 263849 191158 264649
rect 193402 263849 193458 264649
rect 195702 263849 195758 264649
rect 197910 263849 197966 264649
rect 200210 263849 200266 264649
rect 202418 263849 202474 264649
rect 204718 263849 204774 264649
rect 207018 263849 207074 264649
rect 209226 263849 209282 264649
rect 211526 263849 211582 264649
rect 213734 263849 213790 264649
rect 216034 263849 216090 264649
rect 218334 263849 218390 264649
rect 220542 263849 220598 264649
rect 222842 263849 222898 264649
rect 225050 263849 225106 264649
rect 227350 263849 227406 264649
rect 229650 263849 229706 264649
rect 231858 263849 231914 264649
rect 234158 263849 234214 264649
rect 236366 263849 236422 264649
rect 238666 263849 238722 264649
rect 240966 263849 241022 264649
rect 243174 263849 243230 264649
rect 245474 263849 245530 264649
rect 247682 263849 247738 264649
rect 249982 263849 250038 264649
rect 252282 263849 252338 264649
rect 254490 263849 254546 264649
rect 256790 263849 256846 264649
rect 258998 263849 259054 264649
rect 261298 263849 261354 264649
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3330 0 3386 800
rect 3882 0 3938 800
rect 4434 0 4490 800
rect 4986 0 5042 800
rect 5538 0 5594 800
rect 6090 0 6146 800
rect 6550 0 6606 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8206 0 8262 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12990 0 13046 800
rect 13542 0 13598 800
rect 14094 0 14150 800
rect 14646 0 14702 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17314 0 17370 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19430 0 19486 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22650 0 22706 800
rect 23202 0 23258 800
rect 23754 0 23810 800
rect 24306 0 24362 800
rect 24766 0 24822 800
rect 25318 0 25374 800
rect 25870 0 25926 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30654 0 30710 800
rect 31206 0 31262 800
rect 31758 0 31814 800
rect 32310 0 32366 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33874 0 33930 800
rect 34426 0 34482 800
rect 34978 0 35034 800
rect 35530 0 35586 800
rect 36082 0 36138 800
rect 36542 0 36598 800
rect 37094 0 37150 800
rect 37646 0 37702 800
rect 38198 0 38254 800
rect 38750 0 38806 800
rect 39302 0 39358 800
rect 39762 0 39818 800
rect 40314 0 40370 800
rect 40866 0 40922 800
rect 41418 0 41474 800
rect 41970 0 42026 800
rect 42430 0 42486 800
rect 42982 0 43038 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44638 0 44694 800
rect 45190 0 45246 800
rect 45650 0 45706 800
rect 46202 0 46258 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47858 0 47914 800
rect 48410 0 48466 800
rect 48870 0 48926 800
rect 49422 0 49478 800
rect 49974 0 50030 800
rect 50526 0 50582 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 52090 0 52146 800
rect 52642 0 52698 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55310 0 55366 800
rect 55862 0 55918 800
rect 56414 0 56470 800
rect 56966 0 57022 800
rect 57518 0 57574 800
rect 57978 0 58034 800
rect 58530 0 58586 800
rect 59082 0 59138 800
rect 59634 0 59690 800
rect 60186 0 60242 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63406 0 63462 800
rect 63866 0 63922 800
rect 64418 0 64474 800
rect 64970 0 65026 800
rect 65522 0 65578 800
rect 66074 0 66130 800
rect 66534 0 66590 800
rect 67086 0 67142 800
rect 67638 0 67694 800
rect 68190 0 68246 800
rect 68742 0 68798 800
rect 69294 0 69350 800
rect 69754 0 69810 800
rect 70306 0 70362 800
rect 70858 0 70914 800
rect 71410 0 71466 800
rect 71962 0 72018 800
rect 72514 0 72570 800
rect 72974 0 73030 800
rect 73526 0 73582 800
rect 74078 0 74134 800
rect 74630 0 74686 800
rect 75182 0 75238 800
rect 75642 0 75698 800
rect 76194 0 76250 800
rect 76746 0 76802 800
rect 77298 0 77354 800
rect 77850 0 77906 800
rect 78402 0 78458 800
rect 78862 0 78918 800
rect 79414 0 79470 800
rect 79966 0 80022 800
rect 80518 0 80574 800
rect 81070 0 81126 800
rect 81622 0 81678 800
rect 82082 0 82138 800
rect 82634 0 82690 800
rect 83186 0 83242 800
rect 83738 0 83794 800
rect 84290 0 84346 800
rect 84750 0 84806 800
rect 85302 0 85358 800
rect 85854 0 85910 800
rect 86406 0 86462 800
rect 86958 0 87014 800
rect 87510 0 87566 800
rect 87970 0 88026 800
rect 88522 0 88578 800
rect 89074 0 89130 800
rect 89626 0 89682 800
rect 90178 0 90234 800
rect 90638 0 90694 800
rect 91190 0 91246 800
rect 91742 0 91798 800
rect 92294 0 92350 800
rect 92846 0 92902 800
rect 93398 0 93454 800
rect 93858 0 93914 800
rect 94410 0 94466 800
rect 94962 0 95018 800
rect 95514 0 95570 800
rect 96066 0 96122 800
rect 96618 0 96674 800
rect 97078 0 97134 800
rect 97630 0 97686 800
rect 98182 0 98238 800
rect 98734 0 98790 800
rect 99286 0 99342 800
rect 99746 0 99802 800
rect 100298 0 100354 800
rect 100850 0 100906 800
rect 101402 0 101458 800
rect 101954 0 102010 800
rect 102506 0 102562 800
rect 102966 0 103022 800
rect 103518 0 103574 800
rect 104070 0 104126 800
rect 104622 0 104678 800
rect 105174 0 105230 800
rect 105726 0 105782 800
rect 106186 0 106242 800
rect 106738 0 106794 800
rect 107290 0 107346 800
rect 107842 0 107898 800
rect 108394 0 108450 800
rect 108854 0 108910 800
rect 109406 0 109462 800
rect 109958 0 110014 800
rect 110510 0 110566 800
rect 111062 0 111118 800
rect 111614 0 111670 800
rect 112074 0 112130 800
rect 112626 0 112682 800
rect 113178 0 113234 800
rect 113730 0 113786 800
rect 114282 0 114338 800
rect 114834 0 114890 800
rect 115294 0 115350 800
rect 115846 0 115902 800
rect 116398 0 116454 800
rect 116950 0 117006 800
rect 117502 0 117558 800
rect 117962 0 118018 800
rect 118514 0 118570 800
rect 119066 0 119122 800
rect 119618 0 119674 800
rect 120170 0 120226 800
rect 120722 0 120778 800
rect 121182 0 121238 800
rect 121734 0 121790 800
rect 122286 0 122342 800
rect 122838 0 122894 800
rect 123390 0 123446 800
rect 123850 0 123906 800
rect 124402 0 124458 800
rect 124954 0 125010 800
rect 125506 0 125562 800
rect 126058 0 126114 800
rect 126610 0 126666 800
rect 127070 0 127126 800
rect 127622 0 127678 800
rect 128174 0 128230 800
rect 128726 0 128782 800
rect 129278 0 129334 800
rect 129830 0 129886 800
rect 130290 0 130346 800
rect 130842 0 130898 800
rect 131394 0 131450 800
rect 131946 0 132002 800
rect 132498 0 132554 800
rect 132958 0 133014 800
rect 133510 0 133566 800
rect 134062 0 134118 800
rect 134614 0 134670 800
rect 135166 0 135222 800
rect 135718 0 135774 800
rect 136178 0 136234 800
rect 136730 0 136786 800
rect 137282 0 137338 800
rect 137834 0 137890 800
rect 138386 0 138442 800
rect 138938 0 138994 800
rect 139398 0 139454 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 141054 0 141110 800
rect 141606 0 141662 800
rect 142066 0 142122 800
rect 142618 0 142674 800
rect 143170 0 143226 800
rect 143722 0 143778 800
rect 144274 0 144330 800
rect 144826 0 144882 800
rect 145286 0 145342 800
rect 145838 0 145894 800
rect 146390 0 146446 800
rect 146942 0 146998 800
rect 147494 0 147550 800
rect 147954 0 148010 800
rect 148506 0 148562 800
rect 149058 0 149114 800
rect 149610 0 149666 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151174 0 151230 800
rect 151726 0 151782 800
rect 152278 0 152334 800
rect 152830 0 152886 800
rect 153382 0 153438 800
rect 153934 0 153990 800
rect 154394 0 154450 800
rect 154946 0 155002 800
rect 155498 0 155554 800
rect 156050 0 156106 800
rect 156602 0 156658 800
rect 157062 0 157118 800
rect 157614 0 157670 800
rect 158166 0 158222 800
rect 158718 0 158774 800
rect 159270 0 159326 800
rect 159822 0 159878 800
rect 160282 0 160338 800
rect 160834 0 160890 800
rect 161386 0 161442 800
rect 161938 0 161994 800
rect 162490 0 162546 800
rect 163042 0 163098 800
rect 163502 0 163558 800
rect 164054 0 164110 800
rect 164606 0 164662 800
rect 165158 0 165214 800
rect 165710 0 165766 800
rect 166170 0 166226 800
rect 166722 0 166778 800
rect 167274 0 167330 800
rect 167826 0 167882 800
rect 168378 0 168434 800
rect 168930 0 168986 800
rect 169390 0 169446 800
rect 169942 0 169998 800
rect 170494 0 170550 800
rect 171046 0 171102 800
rect 171598 0 171654 800
rect 172150 0 172206 800
rect 172610 0 172666 800
rect 173162 0 173218 800
rect 173714 0 173770 800
rect 174266 0 174322 800
rect 174818 0 174874 800
rect 175278 0 175334 800
rect 175830 0 175886 800
rect 176382 0 176438 800
rect 176934 0 176990 800
rect 177486 0 177542 800
rect 178038 0 178094 800
rect 178498 0 178554 800
rect 179050 0 179106 800
rect 179602 0 179658 800
rect 180154 0 180210 800
rect 180706 0 180762 800
rect 181166 0 181222 800
rect 181718 0 181774 800
rect 182270 0 182326 800
rect 182822 0 182878 800
rect 183374 0 183430 800
rect 183926 0 183982 800
rect 184386 0 184442 800
rect 184938 0 184994 800
rect 185490 0 185546 800
rect 186042 0 186098 800
rect 186594 0 186650 800
rect 187146 0 187202 800
rect 187606 0 187662 800
rect 188158 0 188214 800
rect 188710 0 188766 800
rect 189262 0 189318 800
rect 189814 0 189870 800
rect 190274 0 190330 800
rect 190826 0 190882 800
rect 191378 0 191434 800
rect 191930 0 191986 800
rect 192482 0 192538 800
rect 193034 0 193090 800
rect 193494 0 193550 800
rect 194046 0 194102 800
rect 194598 0 194654 800
rect 195150 0 195206 800
rect 195702 0 195758 800
rect 196254 0 196310 800
rect 196714 0 196770 800
rect 197266 0 197322 800
rect 197818 0 197874 800
rect 198370 0 198426 800
rect 198922 0 198978 800
rect 199382 0 199438 800
rect 199934 0 199990 800
rect 200486 0 200542 800
rect 201038 0 201094 800
rect 201590 0 201646 800
rect 202142 0 202198 800
rect 202602 0 202658 800
rect 203154 0 203210 800
rect 203706 0 203762 800
rect 204258 0 204314 800
rect 204810 0 204866 800
rect 205270 0 205326 800
rect 205822 0 205878 800
rect 206374 0 206430 800
rect 206926 0 206982 800
rect 207478 0 207534 800
rect 208030 0 208086 800
rect 208490 0 208546 800
rect 209042 0 209098 800
rect 209594 0 209650 800
rect 210146 0 210202 800
rect 210698 0 210754 800
rect 211250 0 211306 800
rect 211710 0 211766 800
rect 212262 0 212318 800
rect 212814 0 212870 800
rect 213366 0 213422 800
rect 213918 0 213974 800
rect 214378 0 214434 800
rect 214930 0 214986 800
rect 215482 0 215538 800
rect 216034 0 216090 800
rect 216586 0 216642 800
rect 217138 0 217194 800
rect 217598 0 217654 800
rect 218150 0 218206 800
rect 218702 0 218758 800
rect 219254 0 219310 800
rect 219806 0 219862 800
rect 220358 0 220414 800
rect 220818 0 220874 800
rect 221370 0 221426 800
rect 221922 0 221978 800
rect 222474 0 222530 800
rect 223026 0 223082 800
rect 223486 0 223542 800
rect 224038 0 224094 800
rect 224590 0 224646 800
rect 225142 0 225198 800
rect 225694 0 225750 800
rect 226246 0 226302 800
rect 226706 0 226762 800
rect 227258 0 227314 800
rect 227810 0 227866 800
rect 228362 0 228418 800
rect 228914 0 228970 800
rect 229466 0 229522 800
rect 229926 0 229982 800
rect 230478 0 230534 800
rect 231030 0 231086 800
rect 231582 0 231638 800
rect 232134 0 232190 800
rect 232594 0 232650 800
rect 233146 0 233202 800
rect 233698 0 233754 800
rect 234250 0 234306 800
rect 234802 0 234858 800
rect 235354 0 235410 800
rect 235814 0 235870 800
rect 236366 0 236422 800
rect 236918 0 236974 800
rect 237470 0 237526 800
rect 238022 0 238078 800
rect 238482 0 238538 800
rect 239034 0 239090 800
rect 239586 0 239642 800
rect 240138 0 240194 800
rect 240690 0 240746 800
rect 241242 0 241298 800
rect 241702 0 241758 800
rect 242254 0 242310 800
rect 242806 0 242862 800
rect 243358 0 243414 800
rect 243910 0 243966 800
rect 244462 0 244518 800
rect 244922 0 244978 800
rect 245474 0 245530 800
rect 246026 0 246082 800
rect 246578 0 246634 800
rect 247130 0 247186 800
rect 247590 0 247646 800
rect 248142 0 248198 800
rect 248694 0 248750 800
rect 249246 0 249302 800
rect 249798 0 249854 800
rect 250350 0 250406 800
rect 250810 0 250866 800
rect 251362 0 251418 800
rect 251914 0 251970 800
rect 252466 0 252522 800
rect 253018 0 253074 800
rect 253570 0 253626 800
rect 254030 0 254086 800
rect 254582 0 254638 800
rect 255134 0 255190 800
rect 255686 0 255742 800
rect 256238 0 256294 800
rect 256698 0 256754 800
rect 257250 0 257306 800
rect 257802 0 257858 800
rect 258354 0 258410 800
rect 258906 0 258962 800
rect 259458 0 259514 800
rect 259918 0 259974 800
rect 260470 0 260526 800
rect 261022 0 261078 800
rect 261574 0 261630 800
rect 262126 0 262182 800
<< obsm2 >>
rect 204 263793 1066 263849
rect 1234 263793 3274 263849
rect 3442 263793 5574 263849
rect 5742 263793 7782 263849
rect 7950 263793 10082 263849
rect 10250 263793 12290 263849
rect 12458 263793 14590 263849
rect 14758 263793 16890 263849
rect 17058 263793 19098 263849
rect 19266 263793 21398 263849
rect 21566 263793 23606 263849
rect 23774 263793 25906 263849
rect 26074 263793 28206 263849
rect 28374 263793 30414 263849
rect 30582 263793 32714 263849
rect 32882 263793 34922 263849
rect 35090 263793 37222 263849
rect 37390 263793 39522 263849
rect 39690 263793 41730 263849
rect 41898 263793 44030 263849
rect 44198 263793 46238 263849
rect 46406 263793 48538 263849
rect 48706 263793 50838 263849
rect 51006 263793 53046 263849
rect 53214 263793 55346 263849
rect 55514 263793 57554 263849
rect 57722 263793 59854 263849
rect 60022 263793 62154 263849
rect 62322 263793 64362 263849
rect 64530 263793 66662 263849
rect 66830 263793 68870 263849
rect 69038 263793 71170 263849
rect 71338 263793 73470 263849
rect 73638 263793 75678 263849
rect 75846 263793 77978 263849
rect 78146 263793 80186 263849
rect 80354 263793 82486 263849
rect 82654 263793 84786 263849
rect 84954 263793 86994 263849
rect 87162 263793 89294 263849
rect 89462 263793 91502 263849
rect 91670 263793 93802 263849
rect 93970 263793 96010 263849
rect 96178 263793 98310 263849
rect 98478 263793 100610 263849
rect 100778 263793 102818 263849
rect 102986 263793 105118 263849
rect 105286 263793 107326 263849
rect 107494 263793 109626 263849
rect 109794 263793 111926 263849
rect 112094 263793 114134 263849
rect 114302 263793 116434 263849
rect 116602 263793 118642 263849
rect 118810 263793 120942 263849
rect 121110 263793 123242 263849
rect 123410 263793 125450 263849
rect 125618 263793 127750 263849
rect 127918 263793 129958 263849
rect 130126 263793 132258 263849
rect 132426 263793 134558 263849
rect 134726 263793 136766 263849
rect 136934 263793 139066 263849
rect 139234 263793 141274 263849
rect 141442 263793 143574 263849
rect 143742 263793 145874 263849
rect 146042 263793 148082 263849
rect 148250 263793 150382 263849
rect 150550 263793 152590 263849
rect 152758 263793 154890 263849
rect 155058 263793 157190 263849
rect 157358 263793 159398 263849
rect 159566 263793 161698 263849
rect 161866 263793 163906 263849
rect 164074 263793 166206 263849
rect 166374 263793 168506 263849
rect 168674 263793 170714 263849
rect 170882 263793 173014 263849
rect 173182 263793 175222 263849
rect 175390 263793 177522 263849
rect 177690 263793 179730 263849
rect 179898 263793 182030 263849
rect 182198 263793 184330 263849
rect 184498 263793 186538 263849
rect 186706 263793 188838 263849
rect 189006 263793 191046 263849
rect 191214 263793 193346 263849
rect 193514 263793 195646 263849
rect 195814 263793 197854 263849
rect 198022 263793 200154 263849
rect 200322 263793 202362 263849
rect 202530 263793 204662 263849
rect 204830 263793 206962 263849
rect 207130 263793 209170 263849
rect 209338 263793 211470 263849
rect 211638 263793 213678 263849
rect 213846 263793 215978 263849
rect 216146 263793 218278 263849
rect 218446 263793 220486 263849
rect 220654 263793 222786 263849
rect 222954 263793 224994 263849
rect 225162 263793 227294 263849
rect 227462 263793 229594 263849
rect 229762 263793 231802 263849
rect 231970 263793 234102 263849
rect 234270 263793 236310 263849
rect 236478 263793 238610 263849
rect 238778 263793 240910 263849
rect 241078 263793 243118 263849
rect 243286 263793 245418 263849
rect 245586 263793 247626 263849
rect 247794 263793 249926 263849
rect 250094 263793 252226 263849
rect 252394 263793 254434 263849
rect 254602 263793 256734 263849
rect 256902 263793 258942 263849
rect 259110 263793 261242 263849
rect 261410 263793 262180 263849
rect 204 856 262180 263793
rect 314 800 606 856
rect 774 800 1158 856
rect 1326 800 1710 856
rect 1878 800 2262 856
rect 2430 800 2814 856
rect 2982 800 3274 856
rect 3442 800 3826 856
rect 3994 800 4378 856
rect 4546 800 4930 856
rect 5098 800 5482 856
rect 5650 800 6034 856
rect 6202 800 6494 856
rect 6662 800 7046 856
rect 7214 800 7598 856
rect 7766 800 8150 856
rect 8318 800 8702 856
rect 8870 800 9162 856
rect 9330 800 9714 856
rect 9882 800 10266 856
rect 10434 800 10818 856
rect 10986 800 11370 856
rect 11538 800 11922 856
rect 12090 800 12382 856
rect 12550 800 12934 856
rect 13102 800 13486 856
rect 13654 800 14038 856
rect 14206 800 14590 856
rect 14758 800 15142 856
rect 15310 800 15602 856
rect 15770 800 16154 856
rect 16322 800 16706 856
rect 16874 800 17258 856
rect 17426 800 17810 856
rect 17978 800 18270 856
rect 18438 800 18822 856
rect 18990 800 19374 856
rect 19542 800 19926 856
rect 20094 800 20478 856
rect 20646 800 21030 856
rect 21198 800 21490 856
rect 21658 800 22042 856
rect 22210 800 22594 856
rect 22762 800 23146 856
rect 23314 800 23698 856
rect 23866 800 24250 856
rect 24418 800 24710 856
rect 24878 800 25262 856
rect 25430 800 25814 856
rect 25982 800 26366 856
rect 26534 800 26918 856
rect 27086 800 27378 856
rect 27546 800 27930 856
rect 28098 800 28482 856
rect 28650 800 29034 856
rect 29202 800 29586 856
rect 29754 800 30138 856
rect 30306 800 30598 856
rect 30766 800 31150 856
rect 31318 800 31702 856
rect 31870 800 32254 856
rect 32422 800 32806 856
rect 32974 800 33266 856
rect 33434 800 33818 856
rect 33986 800 34370 856
rect 34538 800 34922 856
rect 35090 800 35474 856
rect 35642 800 36026 856
rect 36194 800 36486 856
rect 36654 800 37038 856
rect 37206 800 37590 856
rect 37758 800 38142 856
rect 38310 800 38694 856
rect 38862 800 39246 856
rect 39414 800 39706 856
rect 39874 800 40258 856
rect 40426 800 40810 856
rect 40978 800 41362 856
rect 41530 800 41914 856
rect 42082 800 42374 856
rect 42542 800 42926 856
rect 43094 800 43478 856
rect 43646 800 44030 856
rect 44198 800 44582 856
rect 44750 800 45134 856
rect 45302 800 45594 856
rect 45762 800 46146 856
rect 46314 800 46698 856
rect 46866 800 47250 856
rect 47418 800 47802 856
rect 47970 800 48354 856
rect 48522 800 48814 856
rect 48982 800 49366 856
rect 49534 800 49918 856
rect 50086 800 50470 856
rect 50638 800 51022 856
rect 51190 800 51482 856
rect 51650 800 52034 856
rect 52202 800 52586 856
rect 52754 800 53138 856
rect 53306 800 53690 856
rect 53858 800 54242 856
rect 54410 800 54702 856
rect 54870 800 55254 856
rect 55422 800 55806 856
rect 55974 800 56358 856
rect 56526 800 56910 856
rect 57078 800 57462 856
rect 57630 800 57922 856
rect 58090 800 58474 856
rect 58642 800 59026 856
rect 59194 800 59578 856
rect 59746 800 60130 856
rect 60298 800 60590 856
rect 60758 800 61142 856
rect 61310 800 61694 856
rect 61862 800 62246 856
rect 62414 800 62798 856
rect 62966 800 63350 856
rect 63518 800 63810 856
rect 63978 800 64362 856
rect 64530 800 64914 856
rect 65082 800 65466 856
rect 65634 800 66018 856
rect 66186 800 66478 856
rect 66646 800 67030 856
rect 67198 800 67582 856
rect 67750 800 68134 856
rect 68302 800 68686 856
rect 68854 800 69238 856
rect 69406 800 69698 856
rect 69866 800 70250 856
rect 70418 800 70802 856
rect 70970 800 71354 856
rect 71522 800 71906 856
rect 72074 800 72458 856
rect 72626 800 72918 856
rect 73086 800 73470 856
rect 73638 800 74022 856
rect 74190 800 74574 856
rect 74742 800 75126 856
rect 75294 800 75586 856
rect 75754 800 76138 856
rect 76306 800 76690 856
rect 76858 800 77242 856
rect 77410 800 77794 856
rect 77962 800 78346 856
rect 78514 800 78806 856
rect 78974 800 79358 856
rect 79526 800 79910 856
rect 80078 800 80462 856
rect 80630 800 81014 856
rect 81182 800 81566 856
rect 81734 800 82026 856
rect 82194 800 82578 856
rect 82746 800 83130 856
rect 83298 800 83682 856
rect 83850 800 84234 856
rect 84402 800 84694 856
rect 84862 800 85246 856
rect 85414 800 85798 856
rect 85966 800 86350 856
rect 86518 800 86902 856
rect 87070 800 87454 856
rect 87622 800 87914 856
rect 88082 800 88466 856
rect 88634 800 89018 856
rect 89186 800 89570 856
rect 89738 800 90122 856
rect 90290 800 90582 856
rect 90750 800 91134 856
rect 91302 800 91686 856
rect 91854 800 92238 856
rect 92406 800 92790 856
rect 92958 800 93342 856
rect 93510 800 93802 856
rect 93970 800 94354 856
rect 94522 800 94906 856
rect 95074 800 95458 856
rect 95626 800 96010 856
rect 96178 800 96562 856
rect 96730 800 97022 856
rect 97190 800 97574 856
rect 97742 800 98126 856
rect 98294 800 98678 856
rect 98846 800 99230 856
rect 99398 800 99690 856
rect 99858 800 100242 856
rect 100410 800 100794 856
rect 100962 800 101346 856
rect 101514 800 101898 856
rect 102066 800 102450 856
rect 102618 800 102910 856
rect 103078 800 103462 856
rect 103630 800 104014 856
rect 104182 800 104566 856
rect 104734 800 105118 856
rect 105286 800 105670 856
rect 105838 800 106130 856
rect 106298 800 106682 856
rect 106850 800 107234 856
rect 107402 800 107786 856
rect 107954 800 108338 856
rect 108506 800 108798 856
rect 108966 800 109350 856
rect 109518 800 109902 856
rect 110070 800 110454 856
rect 110622 800 111006 856
rect 111174 800 111558 856
rect 111726 800 112018 856
rect 112186 800 112570 856
rect 112738 800 113122 856
rect 113290 800 113674 856
rect 113842 800 114226 856
rect 114394 800 114778 856
rect 114946 800 115238 856
rect 115406 800 115790 856
rect 115958 800 116342 856
rect 116510 800 116894 856
rect 117062 800 117446 856
rect 117614 800 117906 856
rect 118074 800 118458 856
rect 118626 800 119010 856
rect 119178 800 119562 856
rect 119730 800 120114 856
rect 120282 800 120666 856
rect 120834 800 121126 856
rect 121294 800 121678 856
rect 121846 800 122230 856
rect 122398 800 122782 856
rect 122950 800 123334 856
rect 123502 800 123794 856
rect 123962 800 124346 856
rect 124514 800 124898 856
rect 125066 800 125450 856
rect 125618 800 126002 856
rect 126170 800 126554 856
rect 126722 800 127014 856
rect 127182 800 127566 856
rect 127734 800 128118 856
rect 128286 800 128670 856
rect 128838 800 129222 856
rect 129390 800 129774 856
rect 129942 800 130234 856
rect 130402 800 130786 856
rect 130954 800 131338 856
rect 131506 800 131890 856
rect 132058 800 132442 856
rect 132610 800 132902 856
rect 133070 800 133454 856
rect 133622 800 134006 856
rect 134174 800 134558 856
rect 134726 800 135110 856
rect 135278 800 135662 856
rect 135830 800 136122 856
rect 136290 800 136674 856
rect 136842 800 137226 856
rect 137394 800 137778 856
rect 137946 800 138330 856
rect 138498 800 138882 856
rect 139050 800 139342 856
rect 139510 800 139894 856
rect 140062 800 140446 856
rect 140614 800 140998 856
rect 141166 800 141550 856
rect 141718 800 142010 856
rect 142178 800 142562 856
rect 142730 800 143114 856
rect 143282 800 143666 856
rect 143834 800 144218 856
rect 144386 800 144770 856
rect 144938 800 145230 856
rect 145398 800 145782 856
rect 145950 800 146334 856
rect 146502 800 146886 856
rect 147054 800 147438 856
rect 147606 800 147898 856
rect 148066 800 148450 856
rect 148618 800 149002 856
rect 149170 800 149554 856
rect 149722 800 150106 856
rect 150274 800 150658 856
rect 150826 800 151118 856
rect 151286 800 151670 856
rect 151838 800 152222 856
rect 152390 800 152774 856
rect 152942 800 153326 856
rect 153494 800 153878 856
rect 154046 800 154338 856
rect 154506 800 154890 856
rect 155058 800 155442 856
rect 155610 800 155994 856
rect 156162 800 156546 856
rect 156714 800 157006 856
rect 157174 800 157558 856
rect 157726 800 158110 856
rect 158278 800 158662 856
rect 158830 800 159214 856
rect 159382 800 159766 856
rect 159934 800 160226 856
rect 160394 800 160778 856
rect 160946 800 161330 856
rect 161498 800 161882 856
rect 162050 800 162434 856
rect 162602 800 162986 856
rect 163154 800 163446 856
rect 163614 800 163998 856
rect 164166 800 164550 856
rect 164718 800 165102 856
rect 165270 800 165654 856
rect 165822 800 166114 856
rect 166282 800 166666 856
rect 166834 800 167218 856
rect 167386 800 167770 856
rect 167938 800 168322 856
rect 168490 800 168874 856
rect 169042 800 169334 856
rect 169502 800 169886 856
rect 170054 800 170438 856
rect 170606 800 170990 856
rect 171158 800 171542 856
rect 171710 800 172094 856
rect 172262 800 172554 856
rect 172722 800 173106 856
rect 173274 800 173658 856
rect 173826 800 174210 856
rect 174378 800 174762 856
rect 174930 800 175222 856
rect 175390 800 175774 856
rect 175942 800 176326 856
rect 176494 800 176878 856
rect 177046 800 177430 856
rect 177598 800 177982 856
rect 178150 800 178442 856
rect 178610 800 178994 856
rect 179162 800 179546 856
rect 179714 800 180098 856
rect 180266 800 180650 856
rect 180818 800 181110 856
rect 181278 800 181662 856
rect 181830 800 182214 856
rect 182382 800 182766 856
rect 182934 800 183318 856
rect 183486 800 183870 856
rect 184038 800 184330 856
rect 184498 800 184882 856
rect 185050 800 185434 856
rect 185602 800 185986 856
rect 186154 800 186538 856
rect 186706 800 187090 856
rect 187258 800 187550 856
rect 187718 800 188102 856
rect 188270 800 188654 856
rect 188822 800 189206 856
rect 189374 800 189758 856
rect 189926 800 190218 856
rect 190386 800 190770 856
rect 190938 800 191322 856
rect 191490 800 191874 856
rect 192042 800 192426 856
rect 192594 800 192978 856
rect 193146 800 193438 856
rect 193606 800 193990 856
rect 194158 800 194542 856
rect 194710 800 195094 856
rect 195262 800 195646 856
rect 195814 800 196198 856
rect 196366 800 196658 856
rect 196826 800 197210 856
rect 197378 800 197762 856
rect 197930 800 198314 856
rect 198482 800 198866 856
rect 199034 800 199326 856
rect 199494 800 199878 856
rect 200046 800 200430 856
rect 200598 800 200982 856
rect 201150 800 201534 856
rect 201702 800 202086 856
rect 202254 800 202546 856
rect 202714 800 203098 856
rect 203266 800 203650 856
rect 203818 800 204202 856
rect 204370 800 204754 856
rect 204922 800 205214 856
rect 205382 800 205766 856
rect 205934 800 206318 856
rect 206486 800 206870 856
rect 207038 800 207422 856
rect 207590 800 207974 856
rect 208142 800 208434 856
rect 208602 800 208986 856
rect 209154 800 209538 856
rect 209706 800 210090 856
rect 210258 800 210642 856
rect 210810 800 211194 856
rect 211362 800 211654 856
rect 211822 800 212206 856
rect 212374 800 212758 856
rect 212926 800 213310 856
rect 213478 800 213862 856
rect 214030 800 214322 856
rect 214490 800 214874 856
rect 215042 800 215426 856
rect 215594 800 215978 856
rect 216146 800 216530 856
rect 216698 800 217082 856
rect 217250 800 217542 856
rect 217710 800 218094 856
rect 218262 800 218646 856
rect 218814 800 219198 856
rect 219366 800 219750 856
rect 219918 800 220302 856
rect 220470 800 220762 856
rect 220930 800 221314 856
rect 221482 800 221866 856
rect 222034 800 222418 856
rect 222586 800 222970 856
rect 223138 800 223430 856
rect 223598 800 223982 856
rect 224150 800 224534 856
rect 224702 800 225086 856
rect 225254 800 225638 856
rect 225806 800 226190 856
rect 226358 800 226650 856
rect 226818 800 227202 856
rect 227370 800 227754 856
rect 227922 800 228306 856
rect 228474 800 228858 856
rect 229026 800 229410 856
rect 229578 800 229870 856
rect 230038 800 230422 856
rect 230590 800 230974 856
rect 231142 800 231526 856
rect 231694 800 232078 856
rect 232246 800 232538 856
rect 232706 800 233090 856
rect 233258 800 233642 856
rect 233810 800 234194 856
rect 234362 800 234746 856
rect 234914 800 235298 856
rect 235466 800 235758 856
rect 235926 800 236310 856
rect 236478 800 236862 856
rect 237030 800 237414 856
rect 237582 800 237966 856
rect 238134 800 238426 856
rect 238594 800 238978 856
rect 239146 800 239530 856
rect 239698 800 240082 856
rect 240250 800 240634 856
rect 240802 800 241186 856
rect 241354 800 241646 856
rect 241814 800 242198 856
rect 242366 800 242750 856
rect 242918 800 243302 856
rect 243470 800 243854 856
rect 244022 800 244406 856
rect 244574 800 244866 856
rect 245034 800 245418 856
rect 245586 800 245970 856
rect 246138 800 246522 856
rect 246690 800 247074 856
rect 247242 800 247534 856
rect 247702 800 248086 856
rect 248254 800 248638 856
rect 248806 800 249190 856
rect 249358 800 249742 856
rect 249910 800 250294 856
rect 250462 800 250754 856
rect 250922 800 251306 856
rect 251474 800 251858 856
rect 252026 800 252410 856
rect 252578 800 252962 856
rect 253130 800 253514 856
rect 253682 800 253974 856
rect 254142 800 254526 856
rect 254694 800 255078 856
rect 255246 800 255630 856
rect 255798 800 256182 856
rect 256350 800 256642 856
rect 256810 800 257194 856
rect 257362 800 257746 856
rect 257914 800 258298 856
rect 258466 800 258850 856
rect 259018 800 259402 856
rect 259570 800 259862 856
rect 260030 800 260414 856
rect 260582 800 260966 856
rect 261134 800 261518 856
rect 261686 800 262070 856
<< metal3 >>
rect 261705 132336 262505 132456
<< obsm3 >>
rect 3141 132536 261705 262241
rect 3141 132256 261625 132536
rect 3141 2143 261705 132256
<< metal4 >>
rect 4208 2128 4528 262256
rect 4868 2176 5188 262208
rect 5528 2176 5848 262208
rect 6188 2176 6508 262208
rect 19568 2128 19888 262256
rect 20228 2176 20548 262208
rect 20888 2176 21208 262208
rect 21548 2176 21868 262208
rect 34928 2128 35248 262256
rect 35588 2176 35908 262208
rect 36248 2176 36568 262208
rect 36908 2176 37228 262208
rect 50288 2128 50608 262256
rect 50948 2176 51268 262208
rect 51608 2176 51928 262208
rect 52268 2176 52588 262208
rect 65648 2128 65968 262256
rect 66308 2176 66628 262208
rect 66968 2176 67288 262208
rect 67628 2176 67948 262208
rect 81008 2128 81328 262256
rect 81668 2176 81988 262208
rect 82328 2176 82648 262208
rect 82988 2176 83308 262208
rect 96368 2128 96688 262256
rect 97028 2176 97348 262208
rect 97688 2176 98008 262208
rect 98348 2176 98668 262208
rect 111728 2128 112048 262256
rect 112388 2176 112708 262208
rect 113048 2176 113368 262208
rect 113708 2176 114028 262208
rect 127088 2128 127408 262256
rect 127748 2176 128068 262208
rect 128408 2176 128728 262208
rect 129068 2176 129388 262208
rect 142448 2128 142768 262256
rect 143108 2176 143428 262208
rect 143768 2176 144088 262208
rect 144428 2176 144748 262208
rect 157808 2128 158128 262256
rect 158468 2176 158788 262208
rect 159128 2176 159448 262208
rect 159788 2176 160108 262208
rect 173168 2128 173488 262256
rect 173828 2176 174148 262208
rect 174488 2176 174808 262208
rect 175148 2176 175468 262208
rect 188528 2128 188848 262256
rect 189188 2176 189508 262208
rect 189848 2176 190168 262208
rect 190508 2176 190828 262208
rect 203888 2128 204208 262256
rect 204548 2176 204868 262208
rect 205208 2176 205528 262208
rect 205868 2176 206188 262208
rect 219248 2128 219568 262256
rect 219908 2176 220228 262208
rect 220568 2176 220888 262208
rect 221228 2176 221548 262208
rect 234608 2128 234928 262256
rect 235268 2176 235588 262208
rect 235928 2176 236248 262208
rect 236588 2176 236908 262208
rect 249968 2128 250288 262256
rect 250628 2176 250948 262208
rect 251288 2176 251608 262208
rect 251948 2176 252268 262208
<< obsm4 >>
rect 21403 27507 21468 186013
rect 21948 27507 34848 186013
rect 35328 27507 35508 186013
rect 35988 27507 36168 186013
rect 36648 27507 36828 186013
rect 37308 27507 50208 186013
rect 50688 27507 50868 186013
rect 51348 27507 51528 186013
rect 52008 27507 52188 186013
rect 52668 27507 65568 186013
rect 66048 27507 66228 186013
rect 66708 27507 66888 186013
rect 67368 27507 67548 186013
rect 68028 27507 80928 186013
rect 81408 27507 81588 186013
rect 82068 27507 82248 186013
rect 82728 27507 82908 186013
rect 83388 27507 96288 186013
rect 96768 27507 96948 186013
rect 97428 27507 97608 186013
rect 98088 27507 98268 186013
rect 98748 27507 111648 186013
rect 112128 27507 112308 186013
rect 112788 27507 112968 186013
rect 113448 27507 113628 186013
rect 114108 27507 127008 186013
rect 127488 27507 127668 186013
rect 128148 27507 128328 186013
rect 128808 27507 128988 186013
rect 129468 27507 142368 186013
rect 142848 27507 143028 186013
rect 143508 27507 143688 186013
rect 144168 27507 144348 186013
rect 144828 27507 157728 186013
rect 158208 27507 158388 186013
rect 158868 27507 159048 186013
rect 159528 27507 159708 186013
rect 160188 27507 173088 186013
rect 173568 27507 173748 186013
rect 174228 27507 174408 186013
rect 174888 27507 175068 186013
rect 175548 27507 188448 186013
rect 188928 27507 189108 186013
rect 189588 27507 189768 186013
rect 190248 27507 190428 186013
rect 190908 27507 203808 186013
<< labels >>
rlabel metal2 s 1122 263849 1178 264649 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 68926 263849 68982 264649 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 75734 263849 75790 264649 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 82542 263849 82598 264649 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 89350 263849 89406 264649 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 96066 263849 96122 264649 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 102874 263849 102930 264649 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 109682 263849 109738 264649 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 116490 263849 116546 264649 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 123298 263849 123354 264649 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 130014 263849 130070 264649 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7838 263849 7894 264649 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 136822 263849 136878 264649 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 143630 263849 143686 264649 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 150438 263849 150494 264649 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 157246 263849 157302 264649 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 163962 263849 164018 264649 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 170770 263849 170826 264649 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 177578 263849 177634 264649 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 184386 263849 184442 264649 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 191102 263849 191158 264649 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 197910 263849 197966 264649 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14646 263849 14702 264649 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 204718 263849 204774 264649 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 211526 263849 211582 264649 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 218334 263849 218390 264649 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 225050 263849 225106 264649 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 231858 263849 231914 264649 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 238666 263849 238722 264649 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 245474 263849 245530 264649 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 252282 263849 252338 264649 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 21454 263849 21510 264649 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 28262 263849 28318 264649 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 34978 263849 35034 264649 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 41786 263849 41842 264649 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 48594 263849 48650 264649 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 55402 263849 55458 264649 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 62210 263849 62266 264649 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3330 263849 3386 264649 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 71226 263849 71282 264649 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 78034 263849 78090 264649 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 84842 263849 84898 264649 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 91558 263849 91614 264649 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 98366 263849 98422 264649 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 105174 263849 105230 264649 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 111982 263849 112038 264649 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 118698 263849 118754 264649 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 125506 263849 125562 264649 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 132314 263849 132370 264649 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 10138 263849 10194 264649 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 139122 263849 139178 264649 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 145930 263849 145986 264649 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 152646 263849 152702 264649 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 159454 263849 159510 264649 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 166262 263849 166318 264649 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 173070 263849 173126 264649 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 179786 263849 179842 264649 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 186594 263849 186650 264649 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 193402 263849 193458 264649 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 200210 263849 200266 264649 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 16946 263849 17002 264649 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 207018 263849 207074 264649 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 213734 263849 213790 264649 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 220542 263849 220598 264649 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 227350 263849 227406 264649 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 234158 263849 234214 264649 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 240966 263849 241022 264649 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 247682 263849 247738 264649 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 254490 263849 254546 264649 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 23662 263849 23718 264649 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 30470 263849 30526 264649 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 37278 263849 37334 264649 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 44086 263849 44142 264649 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 50894 263849 50950 264649 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 57610 263849 57666 264649 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 64418 263849 64474 264649 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5630 263849 5686 264649 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 73526 263849 73582 264649 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 80242 263849 80298 264649 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 87050 263849 87106 264649 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 93858 263849 93914 264649 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 100666 263849 100722 264649 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 107382 263849 107438 264649 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 114190 263849 114246 264649 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 120998 263849 121054 264649 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 127806 263849 127862 264649 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 134614 263849 134670 264649 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 12346 263849 12402 264649 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 141330 263849 141386 264649 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 148138 263849 148194 264649 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 154946 263849 155002 264649 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 161754 263849 161810 264649 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 168562 263849 168618 264649 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 175278 263849 175334 264649 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 182086 263849 182142 264649 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 188894 263849 188950 264649 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 195702 263849 195758 264649 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 202418 263849 202474 264649 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 19154 263849 19210 264649 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 209226 263849 209282 264649 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 216034 263849 216090 264649 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 222842 263849 222898 264649 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 229650 263849 229706 264649 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 236366 263849 236422 264649 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 243174 263849 243230 264649 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 249982 263849 250038 264649 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 256790 263849 256846 264649 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 25962 263849 26018 264649 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 32770 263849 32826 264649 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 39578 263849 39634 264649 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 46294 263849 46350 264649 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 53102 263849 53158 264649 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 59910 263849 59966 264649 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 66718 263849 66774 264649 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 258998 263849 259054 264649 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 261298 263849 261354 264649 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 261705 132336 262505 132456 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 217598 0 217654 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 219254 0 219310 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 224038 0 224094 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 233698 0 233754 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 235354 0 235410 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 238482 0 238538 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 240138 0 240194 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 244922 0 244978 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 246578 0 246634 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 248142 0 248198 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 249798 0 249854 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 251362 0 251418 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 253018 0 253074 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 254582 0 254638 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 257802 0 257858 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 259458 0 259514 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 261022 0 261078 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 164606 0 164662 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 180706 0 180762 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 196714 0 196770 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 203154 0 203210 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 206374 0 206430 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 212814 0 212870 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 216034 0 216090 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 218150 0 218206 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 219806 0 219862 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 221370 0 221426 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 223026 0 223082 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 224590 0 224646 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 226246 0 226302 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 227810 0 227866 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 229466 0 229522 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 231030 0 231086 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 232594 0 232650 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 237470 0 237526 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 239034 0 239090 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 240690 0 240746 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 242254 0 242310 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 243910 0 243966 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 245474 0 245530 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 247130 0 247186 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 248694 0 248750 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 250350 0 250406 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 251914 0 251970 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 253570 0 253626 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 255134 0 255190 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 256698 0 256754 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 258354 0 258410 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 259918 0 259974 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 261574 0 261630 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 163502 0 163558 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 165158 0 165214 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 166722 0 166778 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 176382 0 176438 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 179602 0 179658 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 181166 0 181222 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 182822 0 182878 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 184386 0 184442 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 186042 0 186098 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 187606 0 187662 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 189262 0 189318 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 192482 0 192538 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 194046 0 194102 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 195702 0 195758 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 197266 0 197322 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 198922 0 198978 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 200486 0 200542 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 203706 0 203762 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 205270 0 205326 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 206926 0 206982 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 208490 0 208546 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 210146 0 210202 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 211710 0 211766 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 213366 0 213422 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 214930 0 214986 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 221922 0 221978 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 223486 0 223542 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 239586 0 239642 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 242806 0 242862 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 244462 0 244518 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 247590 0 247646 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 250810 0 250866 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 255686 0 255742 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 258906 0 258962 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 260470 0 260526 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 186594 0 186650 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 196254 0 196310 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 197818 0 197874 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 199382 0 199438 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 204258 0 204314 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 205822 0 205878 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 209042 0 209098 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 210698 0 210754 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 212262 0 212318 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 215482 0 215538 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 249968 2128 250288 262256 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 262256 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 262256 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 262256 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 262256 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 262256 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 262256 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 262256 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 262256 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 234608 2128 234928 262256 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 262256 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 262256 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 262256 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 262256 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 262256 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 262256 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 262256 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 250628 2176 250948 262208 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 262208 6 vccd2
port 626 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 262208 6 vccd2
port 627 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 262208 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 262208 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 262208 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 262208 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 262208 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 262208 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 235268 2176 235588 262208 6 vssd2
port 634 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 262208 6 vssd2
port 635 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 262208 6 vssd2
port 636 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 262208 6 vssd2
port 637 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 262208 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 262208 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 262208 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 262208 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 251288 2176 251608 262208 6 vdda1
port 642 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 262208 6 vdda1
port 643 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 262208 6 vdda1
port 644 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 262208 6 vdda1
port 645 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 262208 6 vdda1
port 646 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 262208 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 262208 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 262208 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 262208 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 235928 2176 236248 262208 6 vssa1
port 651 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 262208 6 vssa1
port 652 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 262208 6 vssa1
port 653 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 262208 6 vssa1
port 654 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 262208 6 vssa1
port 655 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 262208 6 vssa1
port 656 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 262208 6 vssa1
port 657 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 262208 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 251948 2176 252268 262208 6 vdda2
port 659 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 262208 6 vdda2
port 660 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 262208 6 vdda2
port 661 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 262208 6 vdda2
port 662 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 262208 6 vdda2
port 663 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 262208 6 vdda2
port 664 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 262208 6 vdda2
port 665 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 262208 6 vdda2
port 666 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 262208 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 236588 2176 236908 262208 6 vssa2
port 668 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 262208 6 vssa2
port 669 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 262208 6 vssa2
port 670 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 262208 6 vssa2
port 671 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 262208 6 vssa2
port 672 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 262208 6 vssa2
port 673 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 262208 6 vssa2
port 674 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 262208 6 vssa2
port 675 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 262505 264649
string LEFview TRUE
string GDS_FILE /project/openlane/axi_dma/runs/axi_dma/results/magic/axi_dma.gds
string GDS_END 97187170
string GDS_START 1250256
<< end >>

