magic
tech sky130A
magscale 1 2
timestamp 1623988398
<< obsli1 >>
rect 1104 1309 261372 262225
<< obsm1 >>
rect 198 960 262186 262256
<< metal2 >>
rect 1122 263865 1178 264665
rect 3330 263865 3386 264665
rect 5630 263865 5686 264665
rect 7930 263865 7986 264665
rect 10230 263865 10286 264665
rect 12530 263865 12586 264665
rect 14738 263865 14794 264665
rect 17038 263865 17094 264665
rect 19338 263865 19394 264665
rect 21638 263865 21694 264665
rect 23938 263865 23994 264665
rect 26146 263865 26202 264665
rect 28446 263865 28502 264665
rect 30746 263865 30802 264665
rect 33046 263865 33102 264665
rect 35346 263865 35402 264665
rect 37554 263865 37610 264665
rect 39854 263865 39910 264665
rect 42154 263865 42210 264665
rect 44454 263865 44510 264665
rect 46754 263865 46810 264665
rect 48962 263865 49018 264665
rect 51262 263865 51318 264665
rect 53562 263865 53618 264665
rect 55862 263865 55918 264665
rect 58162 263865 58218 264665
rect 60462 263865 60518 264665
rect 62670 263865 62726 264665
rect 64970 263865 65026 264665
rect 67270 263865 67326 264665
rect 69570 263865 69626 264665
rect 71870 263865 71926 264665
rect 74078 263865 74134 264665
rect 76378 263865 76434 264665
rect 78678 263865 78734 264665
rect 80978 263865 81034 264665
rect 83278 263865 83334 264665
rect 85486 263865 85542 264665
rect 87786 263865 87842 264665
rect 90086 263865 90142 264665
rect 92386 263865 92442 264665
rect 94686 263865 94742 264665
rect 96894 263865 96950 264665
rect 99194 263865 99250 264665
rect 101494 263865 101550 264665
rect 103794 263865 103850 264665
rect 106094 263865 106150 264665
rect 108394 263865 108450 264665
rect 110602 263865 110658 264665
rect 112902 263865 112958 264665
rect 115202 263865 115258 264665
rect 117502 263865 117558 264665
rect 119802 263865 119858 264665
rect 122010 263865 122066 264665
rect 124310 263865 124366 264665
rect 126610 263865 126666 264665
rect 128910 263865 128966 264665
rect 131210 263865 131266 264665
rect 133418 263865 133474 264665
rect 135718 263865 135774 264665
rect 138018 263865 138074 264665
rect 140318 263865 140374 264665
rect 142618 263865 142674 264665
rect 144826 263865 144882 264665
rect 147126 263865 147182 264665
rect 149426 263865 149482 264665
rect 151726 263865 151782 264665
rect 154026 263865 154082 264665
rect 156234 263865 156290 264665
rect 158534 263865 158590 264665
rect 160834 263865 160890 264665
rect 163134 263865 163190 264665
rect 165434 263865 165490 264665
rect 167734 263865 167790 264665
rect 169942 263865 169998 264665
rect 172242 263865 172298 264665
rect 174542 263865 174598 264665
rect 176842 263865 176898 264665
rect 179142 263865 179198 264665
rect 181350 263865 181406 264665
rect 183650 263865 183706 264665
rect 185950 263865 186006 264665
rect 188250 263865 188306 264665
rect 190550 263865 190606 264665
rect 192758 263865 192814 264665
rect 195058 263865 195114 264665
rect 197358 263865 197414 264665
rect 199658 263865 199714 264665
rect 201958 263865 202014 264665
rect 204166 263865 204222 264665
rect 206466 263865 206522 264665
rect 208766 263865 208822 264665
rect 211066 263865 211122 264665
rect 213366 263865 213422 264665
rect 215666 263865 215722 264665
rect 217874 263865 217930 264665
rect 220174 263865 220230 264665
rect 222474 263865 222530 264665
rect 224774 263865 224830 264665
rect 227074 263865 227130 264665
rect 229282 263865 229338 264665
rect 231582 263865 231638 264665
rect 233882 263865 233938 264665
rect 236182 263865 236238 264665
rect 238482 263865 238538 264665
rect 240690 263865 240746 264665
rect 242990 263865 243046 264665
rect 245290 263865 245346 264665
rect 247590 263865 247646 264665
rect 249890 263865 249946 264665
rect 252098 263865 252154 264665
rect 254398 263865 254454 264665
rect 256698 263865 256754 264665
rect 258998 263865 259054 264665
rect 261298 263865 261354 264665
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3330 0 3386 800
rect 3882 0 3938 800
rect 4434 0 4490 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5998 0 6054 800
rect 6550 0 6606 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12438 0 12494 800
rect 12990 0 13046 800
rect 13450 0 13506 800
rect 14002 0 14058 800
rect 14554 0 14610 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18786 0 18842 800
rect 19338 0 19394 800
rect 19890 0 19946 800
rect 20442 0 20498 800
rect 20994 0 21050 800
rect 21454 0 21510 800
rect 22006 0 22062 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23662 0 23718 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26790 0 26846 800
rect 27342 0 27398 800
rect 27894 0 27950 800
rect 28446 0 28502 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 30010 0 30066 800
rect 30562 0 30618 800
rect 31114 0 31170 800
rect 31666 0 31722 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35346 0 35402 800
rect 35898 0 35954 800
rect 36450 0 36506 800
rect 37002 0 37058 800
rect 37462 0 37518 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41234 0 41290 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43350 0 43406 800
rect 43902 0 43958 800
rect 44454 0 44510 800
rect 45006 0 45062 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46570 0 46626 800
rect 47122 0 47178 800
rect 47674 0 47730 800
rect 48134 0 48190 800
rect 48686 0 48742 800
rect 49238 0 49294 800
rect 49790 0 49846 800
rect 50342 0 50398 800
rect 50802 0 50858 800
rect 51354 0 51410 800
rect 51906 0 51962 800
rect 52458 0 52514 800
rect 53010 0 53066 800
rect 53470 0 53526 800
rect 54022 0 54078 800
rect 54574 0 54630 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58806 0 58862 800
rect 59358 0 59414 800
rect 59910 0 59966 800
rect 60462 0 60518 800
rect 61014 0 61070 800
rect 61474 0 61530 800
rect 62026 0 62082 800
rect 62578 0 62634 800
rect 63130 0 63186 800
rect 63682 0 63738 800
rect 64142 0 64198 800
rect 64694 0 64750 800
rect 65246 0 65302 800
rect 65798 0 65854 800
rect 66350 0 66406 800
rect 66810 0 66866 800
rect 67362 0 67418 800
rect 67914 0 67970 800
rect 68466 0 68522 800
rect 69018 0 69074 800
rect 69478 0 69534 800
rect 70030 0 70086 800
rect 70582 0 70638 800
rect 71134 0 71190 800
rect 71686 0 71742 800
rect 72146 0 72202 800
rect 72698 0 72754 800
rect 73250 0 73306 800
rect 73802 0 73858 800
rect 74354 0 74410 800
rect 74814 0 74870 800
rect 75366 0 75422 800
rect 75918 0 75974 800
rect 76470 0 76526 800
rect 77022 0 77078 800
rect 77482 0 77538 800
rect 78034 0 78090 800
rect 78586 0 78642 800
rect 79138 0 79194 800
rect 79690 0 79746 800
rect 80150 0 80206 800
rect 80702 0 80758 800
rect 81254 0 81310 800
rect 81806 0 81862 800
rect 82358 0 82414 800
rect 82818 0 82874 800
rect 83370 0 83426 800
rect 83922 0 83978 800
rect 84474 0 84530 800
rect 85026 0 85082 800
rect 85486 0 85542 800
rect 86038 0 86094 800
rect 86590 0 86646 800
rect 87142 0 87198 800
rect 87694 0 87750 800
rect 88154 0 88210 800
rect 88706 0 88762 800
rect 89258 0 89314 800
rect 89810 0 89866 800
rect 90270 0 90326 800
rect 90822 0 90878 800
rect 91374 0 91430 800
rect 91926 0 91982 800
rect 92478 0 92534 800
rect 92938 0 92994 800
rect 93490 0 93546 800
rect 94042 0 94098 800
rect 94594 0 94650 800
rect 95146 0 95202 800
rect 95606 0 95662 800
rect 96158 0 96214 800
rect 96710 0 96766 800
rect 97262 0 97318 800
rect 97814 0 97870 800
rect 98274 0 98330 800
rect 98826 0 98882 800
rect 99378 0 99434 800
rect 99930 0 99986 800
rect 100482 0 100538 800
rect 100942 0 100998 800
rect 101494 0 101550 800
rect 102046 0 102102 800
rect 102598 0 102654 800
rect 103150 0 103206 800
rect 103610 0 103666 800
rect 104162 0 104218 800
rect 104714 0 104770 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106278 0 106334 800
rect 106830 0 106886 800
rect 107382 0 107438 800
rect 107934 0 107990 800
rect 108486 0 108542 800
rect 108946 0 109002 800
rect 109498 0 109554 800
rect 110050 0 110106 800
rect 110602 0 110658 800
rect 111154 0 111210 800
rect 111614 0 111670 800
rect 112166 0 112222 800
rect 112718 0 112774 800
rect 113270 0 113326 800
rect 113822 0 113878 800
rect 114282 0 114338 800
rect 114834 0 114890 800
rect 115386 0 115442 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 116950 0 117006 800
rect 117502 0 117558 800
rect 118054 0 118110 800
rect 118606 0 118662 800
rect 119158 0 119214 800
rect 119618 0 119674 800
rect 120170 0 120226 800
rect 120722 0 120778 800
rect 121274 0 121330 800
rect 121826 0 121882 800
rect 122286 0 122342 800
rect 122838 0 122894 800
rect 123390 0 123446 800
rect 123942 0 123998 800
rect 124494 0 124550 800
rect 124954 0 125010 800
rect 125506 0 125562 800
rect 126058 0 126114 800
rect 126610 0 126666 800
rect 127162 0 127218 800
rect 127622 0 127678 800
rect 128174 0 128230 800
rect 128726 0 128782 800
rect 129278 0 129334 800
rect 129830 0 129886 800
rect 130290 0 130346 800
rect 130842 0 130898 800
rect 131394 0 131450 800
rect 131946 0 132002 800
rect 132498 0 132554 800
rect 132958 0 133014 800
rect 133510 0 133566 800
rect 134062 0 134118 800
rect 134614 0 134670 800
rect 135166 0 135222 800
rect 135626 0 135682 800
rect 136178 0 136234 800
rect 136730 0 136786 800
rect 137282 0 137338 800
rect 137834 0 137890 800
rect 138294 0 138350 800
rect 138846 0 138902 800
rect 139398 0 139454 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 140962 0 141018 800
rect 141514 0 141570 800
rect 142066 0 142122 800
rect 142618 0 142674 800
rect 143170 0 143226 800
rect 143630 0 143686 800
rect 144182 0 144238 800
rect 144734 0 144790 800
rect 145286 0 145342 800
rect 145838 0 145894 800
rect 146298 0 146354 800
rect 146850 0 146906 800
rect 147402 0 147458 800
rect 147954 0 148010 800
rect 148506 0 148562 800
rect 148966 0 149022 800
rect 149518 0 149574 800
rect 150070 0 150126 800
rect 150622 0 150678 800
rect 151174 0 151230 800
rect 151634 0 151690 800
rect 152186 0 152242 800
rect 152738 0 152794 800
rect 153290 0 153346 800
rect 153842 0 153898 800
rect 154302 0 154358 800
rect 154854 0 154910 800
rect 155406 0 155462 800
rect 155958 0 156014 800
rect 156510 0 156566 800
rect 156970 0 157026 800
rect 157522 0 157578 800
rect 158074 0 158130 800
rect 158626 0 158682 800
rect 159178 0 159234 800
rect 159638 0 159694 800
rect 160190 0 160246 800
rect 160742 0 160798 800
rect 161294 0 161350 800
rect 161846 0 161902 800
rect 162306 0 162362 800
rect 162858 0 162914 800
rect 163410 0 163466 800
rect 163962 0 164018 800
rect 164514 0 164570 800
rect 164974 0 165030 800
rect 165526 0 165582 800
rect 166078 0 166134 800
rect 166630 0 166686 800
rect 167182 0 167238 800
rect 167642 0 167698 800
rect 168194 0 168250 800
rect 168746 0 168802 800
rect 169298 0 169354 800
rect 169850 0 169906 800
rect 170310 0 170366 800
rect 170862 0 170918 800
rect 171414 0 171470 800
rect 171966 0 172022 800
rect 172518 0 172574 800
rect 172978 0 173034 800
rect 173530 0 173586 800
rect 174082 0 174138 800
rect 174634 0 174690 800
rect 175186 0 175242 800
rect 175646 0 175702 800
rect 176198 0 176254 800
rect 176750 0 176806 800
rect 177302 0 177358 800
rect 177762 0 177818 800
rect 178314 0 178370 800
rect 178866 0 178922 800
rect 179418 0 179474 800
rect 179970 0 180026 800
rect 180430 0 180486 800
rect 180982 0 181038 800
rect 181534 0 181590 800
rect 182086 0 182142 800
rect 182638 0 182694 800
rect 183098 0 183154 800
rect 183650 0 183706 800
rect 184202 0 184258 800
rect 184754 0 184810 800
rect 185306 0 185362 800
rect 185766 0 185822 800
rect 186318 0 186374 800
rect 186870 0 186926 800
rect 187422 0 187478 800
rect 187974 0 188030 800
rect 188434 0 188490 800
rect 188986 0 189042 800
rect 189538 0 189594 800
rect 190090 0 190146 800
rect 190642 0 190698 800
rect 191102 0 191158 800
rect 191654 0 191710 800
rect 192206 0 192262 800
rect 192758 0 192814 800
rect 193310 0 193366 800
rect 193770 0 193826 800
rect 194322 0 194378 800
rect 194874 0 194930 800
rect 195426 0 195482 800
rect 195978 0 196034 800
rect 196438 0 196494 800
rect 196990 0 197046 800
rect 197542 0 197598 800
rect 198094 0 198150 800
rect 198646 0 198702 800
rect 199106 0 199162 800
rect 199658 0 199714 800
rect 200210 0 200266 800
rect 200762 0 200818 800
rect 201314 0 201370 800
rect 201774 0 201830 800
rect 202326 0 202382 800
rect 202878 0 202934 800
rect 203430 0 203486 800
rect 203982 0 204038 800
rect 204442 0 204498 800
rect 204994 0 205050 800
rect 205546 0 205602 800
rect 206098 0 206154 800
rect 206650 0 206706 800
rect 207110 0 207166 800
rect 207662 0 207718 800
rect 208214 0 208270 800
rect 208766 0 208822 800
rect 209318 0 209374 800
rect 209778 0 209834 800
rect 210330 0 210386 800
rect 210882 0 210938 800
rect 211434 0 211490 800
rect 211986 0 212042 800
rect 212446 0 212502 800
rect 212998 0 213054 800
rect 213550 0 213606 800
rect 214102 0 214158 800
rect 214654 0 214710 800
rect 215114 0 215170 800
rect 215666 0 215722 800
rect 216218 0 216274 800
rect 216770 0 216826 800
rect 217322 0 217378 800
rect 217782 0 217838 800
rect 218334 0 218390 800
rect 218886 0 218942 800
rect 219438 0 219494 800
rect 219990 0 220046 800
rect 220450 0 220506 800
rect 221002 0 221058 800
rect 221554 0 221610 800
rect 222106 0 222162 800
rect 222658 0 222714 800
rect 223118 0 223174 800
rect 223670 0 223726 800
rect 224222 0 224278 800
rect 224774 0 224830 800
rect 225326 0 225382 800
rect 225786 0 225842 800
rect 226338 0 226394 800
rect 226890 0 226946 800
rect 227442 0 227498 800
rect 227994 0 228050 800
rect 228454 0 228510 800
rect 229006 0 229062 800
rect 229558 0 229614 800
rect 230110 0 230166 800
rect 230662 0 230718 800
rect 231122 0 231178 800
rect 231674 0 231730 800
rect 232226 0 232282 800
rect 232778 0 232834 800
rect 233330 0 233386 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234894 0 234950 800
rect 235446 0 235502 800
rect 235998 0 236054 800
rect 236458 0 236514 800
rect 237010 0 237066 800
rect 237562 0 237618 800
rect 238114 0 238170 800
rect 238666 0 238722 800
rect 239126 0 239182 800
rect 239678 0 239734 800
rect 240230 0 240286 800
rect 240782 0 240838 800
rect 241334 0 241390 800
rect 241794 0 241850 800
rect 242346 0 242402 800
rect 242898 0 242954 800
rect 243450 0 243506 800
rect 244002 0 244058 800
rect 244462 0 244518 800
rect 245014 0 245070 800
rect 245566 0 245622 800
rect 246118 0 246174 800
rect 246670 0 246726 800
rect 247130 0 247186 800
rect 247682 0 247738 800
rect 248234 0 248290 800
rect 248786 0 248842 800
rect 249338 0 249394 800
rect 249798 0 249854 800
rect 250350 0 250406 800
rect 250902 0 250958 800
rect 251454 0 251510 800
rect 252006 0 252062 800
rect 252466 0 252522 800
rect 253018 0 253074 800
rect 253570 0 253626 800
rect 254122 0 254178 800
rect 254674 0 254730 800
rect 255134 0 255190 800
rect 255686 0 255742 800
rect 256238 0 256294 800
rect 256790 0 256846 800
rect 257342 0 257398 800
rect 257802 0 257858 800
rect 258354 0 258410 800
rect 258906 0 258962 800
rect 259458 0 259514 800
rect 260010 0 260066 800
rect 260470 0 260526 800
rect 261022 0 261078 800
rect 261574 0 261630 800
rect 262126 0 262182 800
<< obsm2 >>
rect 204 263809 1066 263865
rect 1234 263809 3274 263865
rect 3442 263809 5574 263865
rect 5742 263809 7874 263865
rect 8042 263809 10174 263865
rect 10342 263809 12474 263865
rect 12642 263809 14682 263865
rect 14850 263809 16982 263865
rect 17150 263809 19282 263865
rect 19450 263809 21582 263865
rect 21750 263809 23882 263865
rect 24050 263809 26090 263865
rect 26258 263809 28390 263865
rect 28558 263809 30690 263865
rect 30858 263809 32990 263865
rect 33158 263809 35290 263865
rect 35458 263809 37498 263865
rect 37666 263809 39798 263865
rect 39966 263809 42098 263865
rect 42266 263809 44398 263865
rect 44566 263809 46698 263865
rect 46866 263809 48906 263865
rect 49074 263809 51206 263865
rect 51374 263809 53506 263865
rect 53674 263809 55806 263865
rect 55974 263809 58106 263865
rect 58274 263809 60406 263865
rect 60574 263809 62614 263865
rect 62782 263809 64914 263865
rect 65082 263809 67214 263865
rect 67382 263809 69514 263865
rect 69682 263809 71814 263865
rect 71982 263809 74022 263865
rect 74190 263809 76322 263865
rect 76490 263809 78622 263865
rect 78790 263809 80922 263865
rect 81090 263809 83222 263865
rect 83390 263809 85430 263865
rect 85598 263809 87730 263865
rect 87898 263809 90030 263865
rect 90198 263809 92330 263865
rect 92498 263809 94630 263865
rect 94798 263809 96838 263865
rect 97006 263809 99138 263865
rect 99306 263809 101438 263865
rect 101606 263809 103738 263865
rect 103906 263809 106038 263865
rect 106206 263809 108338 263865
rect 108506 263809 110546 263865
rect 110714 263809 112846 263865
rect 113014 263809 115146 263865
rect 115314 263809 117446 263865
rect 117614 263809 119746 263865
rect 119914 263809 121954 263865
rect 122122 263809 124254 263865
rect 124422 263809 126554 263865
rect 126722 263809 128854 263865
rect 129022 263809 131154 263865
rect 131322 263809 133362 263865
rect 133530 263809 135662 263865
rect 135830 263809 137962 263865
rect 138130 263809 140262 263865
rect 140430 263809 142562 263865
rect 142730 263809 144770 263865
rect 144938 263809 147070 263865
rect 147238 263809 149370 263865
rect 149538 263809 151670 263865
rect 151838 263809 153970 263865
rect 154138 263809 156178 263865
rect 156346 263809 158478 263865
rect 158646 263809 160778 263865
rect 160946 263809 163078 263865
rect 163246 263809 165378 263865
rect 165546 263809 167678 263865
rect 167846 263809 169886 263865
rect 170054 263809 172186 263865
rect 172354 263809 174486 263865
rect 174654 263809 176786 263865
rect 176954 263809 179086 263865
rect 179254 263809 181294 263865
rect 181462 263809 183594 263865
rect 183762 263809 185894 263865
rect 186062 263809 188194 263865
rect 188362 263809 190494 263865
rect 190662 263809 192702 263865
rect 192870 263809 195002 263865
rect 195170 263809 197302 263865
rect 197470 263809 199602 263865
rect 199770 263809 201902 263865
rect 202070 263809 204110 263865
rect 204278 263809 206410 263865
rect 206578 263809 208710 263865
rect 208878 263809 211010 263865
rect 211178 263809 213310 263865
rect 213478 263809 215610 263865
rect 215778 263809 217818 263865
rect 217986 263809 220118 263865
rect 220286 263809 222418 263865
rect 222586 263809 224718 263865
rect 224886 263809 227018 263865
rect 227186 263809 229226 263865
rect 229394 263809 231526 263865
rect 231694 263809 233826 263865
rect 233994 263809 236126 263865
rect 236294 263809 238426 263865
rect 238594 263809 240634 263865
rect 240802 263809 242934 263865
rect 243102 263809 245234 263865
rect 245402 263809 247534 263865
rect 247702 263809 249834 263865
rect 250002 263809 252042 263865
rect 252210 263809 254342 263865
rect 254510 263809 256642 263865
rect 256810 263809 258942 263865
rect 259110 263809 261242 263865
rect 261410 263809 262180 263865
rect 204 856 262180 263809
rect 314 800 606 856
rect 774 800 1158 856
rect 1326 800 1710 856
rect 1878 800 2262 856
rect 2430 800 2722 856
rect 2890 800 3274 856
rect 3442 800 3826 856
rect 3994 800 4378 856
rect 4546 800 4930 856
rect 5098 800 5390 856
rect 5558 800 5942 856
rect 6110 800 6494 856
rect 6662 800 7046 856
rect 7214 800 7598 856
rect 7766 800 8058 856
rect 8226 800 8610 856
rect 8778 800 9162 856
rect 9330 800 9714 856
rect 9882 800 10266 856
rect 10434 800 10726 856
rect 10894 800 11278 856
rect 11446 800 11830 856
rect 11998 800 12382 856
rect 12550 800 12934 856
rect 13102 800 13394 856
rect 13562 800 13946 856
rect 14114 800 14498 856
rect 14666 800 15050 856
rect 15218 800 15602 856
rect 15770 800 16062 856
rect 16230 800 16614 856
rect 16782 800 17166 856
rect 17334 800 17718 856
rect 17886 800 18270 856
rect 18438 800 18730 856
rect 18898 800 19282 856
rect 19450 800 19834 856
rect 20002 800 20386 856
rect 20554 800 20938 856
rect 21106 800 21398 856
rect 21566 800 21950 856
rect 22118 800 22502 856
rect 22670 800 23054 856
rect 23222 800 23606 856
rect 23774 800 24066 856
rect 24234 800 24618 856
rect 24786 800 25170 856
rect 25338 800 25722 856
rect 25890 800 26274 856
rect 26442 800 26734 856
rect 26902 800 27286 856
rect 27454 800 27838 856
rect 28006 800 28390 856
rect 28558 800 28942 856
rect 29110 800 29402 856
rect 29570 800 29954 856
rect 30122 800 30506 856
rect 30674 800 31058 856
rect 31226 800 31610 856
rect 31778 800 32070 856
rect 32238 800 32622 856
rect 32790 800 33174 856
rect 33342 800 33726 856
rect 33894 800 34278 856
rect 34446 800 34738 856
rect 34906 800 35290 856
rect 35458 800 35842 856
rect 36010 800 36394 856
rect 36562 800 36946 856
rect 37114 800 37406 856
rect 37574 800 37958 856
rect 38126 800 38510 856
rect 38678 800 39062 856
rect 39230 800 39614 856
rect 39782 800 40074 856
rect 40242 800 40626 856
rect 40794 800 41178 856
rect 41346 800 41730 856
rect 41898 800 42282 856
rect 42450 800 42742 856
rect 42910 800 43294 856
rect 43462 800 43846 856
rect 44014 800 44398 856
rect 44566 800 44950 856
rect 45118 800 45410 856
rect 45578 800 45962 856
rect 46130 800 46514 856
rect 46682 800 47066 856
rect 47234 800 47618 856
rect 47786 800 48078 856
rect 48246 800 48630 856
rect 48798 800 49182 856
rect 49350 800 49734 856
rect 49902 800 50286 856
rect 50454 800 50746 856
rect 50914 800 51298 856
rect 51466 800 51850 856
rect 52018 800 52402 856
rect 52570 800 52954 856
rect 53122 800 53414 856
rect 53582 800 53966 856
rect 54134 800 54518 856
rect 54686 800 55070 856
rect 55238 800 55622 856
rect 55790 800 56082 856
rect 56250 800 56634 856
rect 56802 800 57186 856
rect 57354 800 57738 856
rect 57906 800 58290 856
rect 58458 800 58750 856
rect 58918 800 59302 856
rect 59470 800 59854 856
rect 60022 800 60406 856
rect 60574 800 60958 856
rect 61126 800 61418 856
rect 61586 800 61970 856
rect 62138 800 62522 856
rect 62690 800 63074 856
rect 63242 800 63626 856
rect 63794 800 64086 856
rect 64254 800 64638 856
rect 64806 800 65190 856
rect 65358 800 65742 856
rect 65910 800 66294 856
rect 66462 800 66754 856
rect 66922 800 67306 856
rect 67474 800 67858 856
rect 68026 800 68410 856
rect 68578 800 68962 856
rect 69130 800 69422 856
rect 69590 800 69974 856
rect 70142 800 70526 856
rect 70694 800 71078 856
rect 71246 800 71630 856
rect 71798 800 72090 856
rect 72258 800 72642 856
rect 72810 800 73194 856
rect 73362 800 73746 856
rect 73914 800 74298 856
rect 74466 800 74758 856
rect 74926 800 75310 856
rect 75478 800 75862 856
rect 76030 800 76414 856
rect 76582 800 76966 856
rect 77134 800 77426 856
rect 77594 800 77978 856
rect 78146 800 78530 856
rect 78698 800 79082 856
rect 79250 800 79634 856
rect 79802 800 80094 856
rect 80262 800 80646 856
rect 80814 800 81198 856
rect 81366 800 81750 856
rect 81918 800 82302 856
rect 82470 800 82762 856
rect 82930 800 83314 856
rect 83482 800 83866 856
rect 84034 800 84418 856
rect 84586 800 84970 856
rect 85138 800 85430 856
rect 85598 800 85982 856
rect 86150 800 86534 856
rect 86702 800 87086 856
rect 87254 800 87638 856
rect 87806 800 88098 856
rect 88266 800 88650 856
rect 88818 800 89202 856
rect 89370 800 89754 856
rect 89922 800 90214 856
rect 90382 800 90766 856
rect 90934 800 91318 856
rect 91486 800 91870 856
rect 92038 800 92422 856
rect 92590 800 92882 856
rect 93050 800 93434 856
rect 93602 800 93986 856
rect 94154 800 94538 856
rect 94706 800 95090 856
rect 95258 800 95550 856
rect 95718 800 96102 856
rect 96270 800 96654 856
rect 96822 800 97206 856
rect 97374 800 97758 856
rect 97926 800 98218 856
rect 98386 800 98770 856
rect 98938 800 99322 856
rect 99490 800 99874 856
rect 100042 800 100426 856
rect 100594 800 100886 856
rect 101054 800 101438 856
rect 101606 800 101990 856
rect 102158 800 102542 856
rect 102710 800 103094 856
rect 103262 800 103554 856
rect 103722 800 104106 856
rect 104274 800 104658 856
rect 104826 800 105210 856
rect 105378 800 105762 856
rect 105930 800 106222 856
rect 106390 800 106774 856
rect 106942 800 107326 856
rect 107494 800 107878 856
rect 108046 800 108430 856
rect 108598 800 108890 856
rect 109058 800 109442 856
rect 109610 800 109994 856
rect 110162 800 110546 856
rect 110714 800 111098 856
rect 111266 800 111558 856
rect 111726 800 112110 856
rect 112278 800 112662 856
rect 112830 800 113214 856
rect 113382 800 113766 856
rect 113934 800 114226 856
rect 114394 800 114778 856
rect 114946 800 115330 856
rect 115498 800 115882 856
rect 116050 800 116434 856
rect 116602 800 116894 856
rect 117062 800 117446 856
rect 117614 800 117998 856
rect 118166 800 118550 856
rect 118718 800 119102 856
rect 119270 800 119562 856
rect 119730 800 120114 856
rect 120282 800 120666 856
rect 120834 800 121218 856
rect 121386 800 121770 856
rect 121938 800 122230 856
rect 122398 800 122782 856
rect 122950 800 123334 856
rect 123502 800 123886 856
rect 124054 800 124438 856
rect 124606 800 124898 856
rect 125066 800 125450 856
rect 125618 800 126002 856
rect 126170 800 126554 856
rect 126722 800 127106 856
rect 127274 800 127566 856
rect 127734 800 128118 856
rect 128286 800 128670 856
rect 128838 800 129222 856
rect 129390 800 129774 856
rect 129942 800 130234 856
rect 130402 800 130786 856
rect 130954 800 131338 856
rect 131506 800 131890 856
rect 132058 800 132442 856
rect 132610 800 132902 856
rect 133070 800 133454 856
rect 133622 800 134006 856
rect 134174 800 134558 856
rect 134726 800 135110 856
rect 135278 800 135570 856
rect 135738 800 136122 856
rect 136290 800 136674 856
rect 136842 800 137226 856
rect 137394 800 137778 856
rect 137946 800 138238 856
rect 138406 800 138790 856
rect 138958 800 139342 856
rect 139510 800 139894 856
rect 140062 800 140446 856
rect 140614 800 140906 856
rect 141074 800 141458 856
rect 141626 800 142010 856
rect 142178 800 142562 856
rect 142730 800 143114 856
rect 143282 800 143574 856
rect 143742 800 144126 856
rect 144294 800 144678 856
rect 144846 800 145230 856
rect 145398 800 145782 856
rect 145950 800 146242 856
rect 146410 800 146794 856
rect 146962 800 147346 856
rect 147514 800 147898 856
rect 148066 800 148450 856
rect 148618 800 148910 856
rect 149078 800 149462 856
rect 149630 800 150014 856
rect 150182 800 150566 856
rect 150734 800 151118 856
rect 151286 800 151578 856
rect 151746 800 152130 856
rect 152298 800 152682 856
rect 152850 800 153234 856
rect 153402 800 153786 856
rect 153954 800 154246 856
rect 154414 800 154798 856
rect 154966 800 155350 856
rect 155518 800 155902 856
rect 156070 800 156454 856
rect 156622 800 156914 856
rect 157082 800 157466 856
rect 157634 800 158018 856
rect 158186 800 158570 856
rect 158738 800 159122 856
rect 159290 800 159582 856
rect 159750 800 160134 856
rect 160302 800 160686 856
rect 160854 800 161238 856
rect 161406 800 161790 856
rect 161958 800 162250 856
rect 162418 800 162802 856
rect 162970 800 163354 856
rect 163522 800 163906 856
rect 164074 800 164458 856
rect 164626 800 164918 856
rect 165086 800 165470 856
rect 165638 800 166022 856
rect 166190 800 166574 856
rect 166742 800 167126 856
rect 167294 800 167586 856
rect 167754 800 168138 856
rect 168306 800 168690 856
rect 168858 800 169242 856
rect 169410 800 169794 856
rect 169962 800 170254 856
rect 170422 800 170806 856
rect 170974 800 171358 856
rect 171526 800 171910 856
rect 172078 800 172462 856
rect 172630 800 172922 856
rect 173090 800 173474 856
rect 173642 800 174026 856
rect 174194 800 174578 856
rect 174746 800 175130 856
rect 175298 800 175590 856
rect 175758 800 176142 856
rect 176310 800 176694 856
rect 176862 800 177246 856
rect 177414 800 177706 856
rect 177874 800 178258 856
rect 178426 800 178810 856
rect 178978 800 179362 856
rect 179530 800 179914 856
rect 180082 800 180374 856
rect 180542 800 180926 856
rect 181094 800 181478 856
rect 181646 800 182030 856
rect 182198 800 182582 856
rect 182750 800 183042 856
rect 183210 800 183594 856
rect 183762 800 184146 856
rect 184314 800 184698 856
rect 184866 800 185250 856
rect 185418 800 185710 856
rect 185878 800 186262 856
rect 186430 800 186814 856
rect 186982 800 187366 856
rect 187534 800 187918 856
rect 188086 800 188378 856
rect 188546 800 188930 856
rect 189098 800 189482 856
rect 189650 800 190034 856
rect 190202 800 190586 856
rect 190754 800 191046 856
rect 191214 800 191598 856
rect 191766 800 192150 856
rect 192318 800 192702 856
rect 192870 800 193254 856
rect 193422 800 193714 856
rect 193882 800 194266 856
rect 194434 800 194818 856
rect 194986 800 195370 856
rect 195538 800 195922 856
rect 196090 800 196382 856
rect 196550 800 196934 856
rect 197102 800 197486 856
rect 197654 800 198038 856
rect 198206 800 198590 856
rect 198758 800 199050 856
rect 199218 800 199602 856
rect 199770 800 200154 856
rect 200322 800 200706 856
rect 200874 800 201258 856
rect 201426 800 201718 856
rect 201886 800 202270 856
rect 202438 800 202822 856
rect 202990 800 203374 856
rect 203542 800 203926 856
rect 204094 800 204386 856
rect 204554 800 204938 856
rect 205106 800 205490 856
rect 205658 800 206042 856
rect 206210 800 206594 856
rect 206762 800 207054 856
rect 207222 800 207606 856
rect 207774 800 208158 856
rect 208326 800 208710 856
rect 208878 800 209262 856
rect 209430 800 209722 856
rect 209890 800 210274 856
rect 210442 800 210826 856
rect 210994 800 211378 856
rect 211546 800 211930 856
rect 212098 800 212390 856
rect 212558 800 212942 856
rect 213110 800 213494 856
rect 213662 800 214046 856
rect 214214 800 214598 856
rect 214766 800 215058 856
rect 215226 800 215610 856
rect 215778 800 216162 856
rect 216330 800 216714 856
rect 216882 800 217266 856
rect 217434 800 217726 856
rect 217894 800 218278 856
rect 218446 800 218830 856
rect 218998 800 219382 856
rect 219550 800 219934 856
rect 220102 800 220394 856
rect 220562 800 220946 856
rect 221114 800 221498 856
rect 221666 800 222050 856
rect 222218 800 222602 856
rect 222770 800 223062 856
rect 223230 800 223614 856
rect 223782 800 224166 856
rect 224334 800 224718 856
rect 224886 800 225270 856
rect 225438 800 225730 856
rect 225898 800 226282 856
rect 226450 800 226834 856
rect 227002 800 227386 856
rect 227554 800 227938 856
rect 228106 800 228398 856
rect 228566 800 228950 856
rect 229118 800 229502 856
rect 229670 800 230054 856
rect 230222 800 230606 856
rect 230774 800 231066 856
rect 231234 800 231618 856
rect 231786 800 232170 856
rect 232338 800 232722 856
rect 232890 800 233274 856
rect 233442 800 233734 856
rect 233902 800 234286 856
rect 234454 800 234838 856
rect 235006 800 235390 856
rect 235558 800 235942 856
rect 236110 800 236402 856
rect 236570 800 236954 856
rect 237122 800 237506 856
rect 237674 800 238058 856
rect 238226 800 238610 856
rect 238778 800 239070 856
rect 239238 800 239622 856
rect 239790 800 240174 856
rect 240342 800 240726 856
rect 240894 800 241278 856
rect 241446 800 241738 856
rect 241906 800 242290 856
rect 242458 800 242842 856
rect 243010 800 243394 856
rect 243562 800 243946 856
rect 244114 800 244406 856
rect 244574 800 244958 856
rect 245126 800 245510 856
rect 245678 800 246062 856
rect 246230 800 246614 856
rect 246782 800 247074 856
rect 247242 800 247626 856
rect 247794 800 248178 856
rect 248346 800 248730 856
rect 248898 800 249282 856
rect 249450 800 249742 856
rect 249910 800 250294 856
rect 250462 800 250846 856
rect 251014 800 251398 856
rect 251566 800 251950 856
rect 252118 800 252410 856
rect 252578 800 252962 856
rect 253130 800 253514 856
rect 253682 800 254066 856
rect 254234 800 254618 856
rect 254786 800 255078 856
rect 255246 800 255630 856
rect 255798 800 256182 856
rect 256350 800 256734 856
rect 256902 800 257286 856
rect 257454 800 257746 856
rect 257914 800 258298 856
rect 258466 800 258850 856
rect 259018 800 259402 856
rect 259570 800 259954 856
rect 260122 800 260414 856
rect 260582 800 260966 856
rect 261134 800 261518 856
rect 261686 800 262070 856
<< obsm3 >>
rect 4208 1395 260071 262241
<< metal4 >>
rect 4208 2128 4528 262256
rect 4868 2176 5188 262208
rect 5528 2176 5848 262208
rect 6188 2176 6508 262208
rect 19568 2128 19888 262256
rect 20228 2176 20548 262208
rect 20888 2176 21208 262208
rect 21548 2176 21868 262208
rect 34928 2128 35248 262256
rect 35588 2176 35908 262208
rect 36248 2176 36568 262208
rect 36908 2176 37228 262208
rect 50288 2128 50608 262256
rect 50948 2176 51268 262208
rect 51608 2176 51928 262208
rect 52268 2176 52588 262208
rect 65648 2128 65968 262256
rect 66308 2176 66628 262208
rect 66968 2176 67288 262208
rect 67628 2176 67948 262208
rect 81008 2128 81328 262256
rect 81668 2176 81988 262208
rect 82328 2176 82648 262208
rect 82988 2176 83308 262208
rect 96368 2128 96688 262256
rect 97028 2176 97348 262208
rect 97688 2176 98008 262208
rect 98348 2176 98668 262208
rect 111728 2128 112048 262256
rect 112388 2176 112708 262208
rect 113048 2176 113368 262208
rect 113708 2176 114028 262208
rect 127088 2128 127408 262256
rect 127748 2176 128068 262208
rect 128408 2176 128728 262208
rect 129068 2176 129388 262208
rect 142448 2128 142768 262256
rect 143108 2176 143428 262208
rect 143768 2176 144088 262208
rect 144428 2176 144748 262208
rect 157808 2128 158128 262256
rect 158468 2176 158788 262208
rect 159128 2176 159448 262208
rect 159788 2176 160108 262208
rect 173168 2128 173488 262256
rect 173828 2176 174148 262208
rect 174488 2176 174808 262208
rect 175148 2176 175468 262208
rect 188528 2128 188848 262256
rect 189188 2176 189508 262208
rect 189848 2176 190168 262208
rect 190508 2176 190828 262208
rect 203888 2128 204208 262256
rect 204548 2176 204868 262208
rect 205208 2176 205528 262208
rect 205868 2176 206188 262208
rect 219248 2128 219568 262256
rect 219908 2176 220228 262208
rect 220568 2176 220888 262208
rect 221228 2176 221548 262208
rect 234608 2128 234928 262256
rect 235268 2176 235588 262208
rect 235928 2176 236248 262208
rect 236588 2176 236908 262208
rect 249968 2128 250288 262256
rect 250628 2176 250948 262208
rect 251288 2176 251608 262208
rect 251948 2176 252268 262208
<< obsm4 >>
rect 19379 18803 19488 245037
rect 19968 18803 20148 245037
rect 20628 18803 20808 245037
rect 21288 18803 21468 245037
rect 21948 18803 34848 245037
rect 35328 18803 35508 245037
rect 35988 18803 36168 245037
rect 36648 18803 36828 245037
rect 37308 18803 50208 245037
rect 50688 18803 50868 245037
rect 51348 18803 51528 245037
rect 52008 18803 52188 245037
rect 52668 18803 65568 245037
rect 66048 18803 66228 245037
rect 66708 18803 66888 245037
rect 67368 18803 67548 245037
rect 68028 18803 80928 245037
rect 81408 18803 81588 245037
rect 82068 18803 82248 245037
rect 82728 18803 82908 245037
rect 83388 18803 96288 245037
rect 96768 18803 96948 245037
rect 97428 18803 97608 245037
rect 98088 18803 98268 245037
rect 98748 18803 111648 245037
rect 112128 18803 112308 245037
rect 112788 18803 112968 245037
rect 113448 18803 113628 245037
rect 114108 18803 127008 245037
rect 127488 18803 127668 245037
rect 128148 18803 128328 245037
rect 128808 18803 128988 245037
rect 129468 18803 142368 245037
rect 142848 18803 143028 245037
rect 143508 18803 143688 245037
rect 144168 18803 144348 245037
rect 144828 18803 157728 245037
rect 158208 18803 158388 245037
rect 158868 18803 159048 245037
rect 159528 18803 159708 245037
rect 160188 18803 173088 245037
rect 173568 18803 173748 245037
rect 174228 18803 174408 245037
rect 174888 18803 175068 245037
rect 175548 18803 188448 245037
rect 188928 18803 189108 245037
rect 189588 18803 189768 245037
rect 190248 18803 190428 245037
rect 190908 18803 203808 245037
rect 204288 18803 204468 245037
rect 204948 18803 205128 245037
rect 205608 18803 205788 245037
rect 206268 18803 219168 245037
rect 219648 18803 219828 245037
rect 220308 18803 220488 245037
rect 220968 18803 221148 245037
rect 221628 18803 222213 245037
<< labels >>
rlabel metal2 s 1122 263865 1178 264665 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 69570 263865 69626 264665 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 76378 263865 76434 264665 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 83278 263865 83334 264665 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 90086 263865 90142 264665 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 96894 263865 96950 264665 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 103794 263865 103850 264665 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 110602 263865 110658 264665 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 117502 263865 117558 264665 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 124310 263865 124366 264665 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 131210 263865 131266 264665 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7930 263865 7986 264665 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 138018 263865 138074 264665 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 144826 263865 144882 264665 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 151726 263865 151782 264665 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 158534 263865 158590 264665 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 165434 263865 165490 264665 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 172242 263865 172298 264665 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 179142 263865 179198 264665 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 185950 263865 186006 264665 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 192758 263865 192814 264665 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 199658 263865 199714 264665 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14738 263865 14794 264665 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 206466 263865 206522 264665 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 213366 263865 213422 264665 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 220174 263865 220230 264665 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 227074 263865 227130 264665 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 233882 263865 233938 264665 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 240690 263865 240746 264665 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 247590 263865 247646 264665 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 254398 263865 254454 264665 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 21638 263865 21694 264665 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 28446 263865 28502 264665 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 35346 263865 35402 264665 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 42154 263865 42210 264665 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 48962 263865 49018 264665 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 55862 263865 55918 264665 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 62670 263865 62726 264665 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3330 263865 3386 264665 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 71870 263865 71926 264665 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 78678 263865 78734 264665 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 85486 263865 85542 264665 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 92386 263865 92442 264665 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 99194 263865 99250 264665 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 106094 263865 106150 264665 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 112902 263865 112958 264665 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 119802 263865 119858 264665 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 126610 263865 126666 264665 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 133418 263865 133474 264665 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 10230 263865 10286 264665 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 140318 263865 140374 264665 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 147126 263865 147182 264665 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 154026 263865 154082 264665 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 160834 263865 160890 264665 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 167734 263865 167790 264665 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 174542 263865 174598 264665 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 181350 263865 181406 264665 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 188250 263865 188306 264665 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 195058 263865 195114 264665 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 201958 263865 202014 264665 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 17038 263865 17094 264665 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 208766 263865 208822 264665 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 215666 263865 215722 264665 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 222474 263865 222530 264665 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 229282 263865 229338 264665 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 236182 263865 236238 264665 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 242990 263865 243046 264665 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 249890 263865 249946 264665 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 256698 263865 256754 264665 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 23938 263865 23994 264665 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 30746 263865 30802 264665 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 37554 263865 37610 264665 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 44454 263865 44510 264665 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 51262 263865 51318 264665 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 58162 263865 58218 264665 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 64970 263865 65026 264665 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5630 263865 5686 264665 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 74078 263865 74134 264665 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 80978 263865 81034 264665 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 87786 263865 87842 264665 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 94686 263865 94742 264665 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 101494 263865 101550 264665 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 108394 263865 108450 264665 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 115202 263865 115258 264665 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 122010 263865 122066 264665 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 128910 263865 128966 264665 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 135718 263865 135774 264665 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 12530 263865 12586 264665 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 142618 263865 142674 264665 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 149426 263865 149482 264665 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 156234 263865 156290 264665 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 163134 263865 163190 264665 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 169942 263865 169998 264665 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 176842 263865 176898 264665 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 183650 263865 183706 264665 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 190550 263865 190606 264665 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 197358 263865 197414 264665 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 204166 263865 204222 264665 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 19338 263865 19394 264665 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 211066 263865 211122 264665 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 217874 263865 217930 264665 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 224774 263865 224830 264665 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 231582 263865 231638 264665 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 238482 263865 238538 264665 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 245290 263865 245346 264665 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 252098 263865 252154 264665 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 258998 263865 259054 264665 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 26146 263865 26202 264665 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 33046 263865 33102 264665 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 39854 263865 39910 264665 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 46754 263865 46810 264665 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 53562 263865 53618 264665 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 60462 263865 60518 264665 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 67270 263865 67326 264665 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 261298 263865 261354 264665 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 261574 0 261630 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 262126 0 262182 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 216770 0 216826 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 219990 0 220046 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 229558 0 229614 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 234342 0 234398 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 235998 0 236054 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 242346 0 242402 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 247130 0 247186 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 248786 0 248842 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 250350 0 250406 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 252006 0 252062 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 253570 0 253626 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 255134 0 255190 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 260010 0 260066 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 179970 0 180026 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 181534 0 181590 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 200762 0 200818 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 202326 0 202382 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 203982 0 204038 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 205546 0 205602 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 207110 0 207166 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 208766 0 208822 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 213550 0 213606 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 217322 0 217378 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 218886 0 218942 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 220450 0 220506 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 222106 0 222162 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 223670 0 223726 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 225326 0 225382 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 226890 0 226946 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 228454 0 228510 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 230110 0 230166 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 231674 0 231730 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 234894 0 234950 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 236458 0 236514 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 238114 0 238170 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 239678 0 239734 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 241334 0 241390 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 242898 0 242954 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 244462 0 244518 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 246118 0 246174 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 247682 0 247738 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 249338 0 249394 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 250902 0 250958 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 252466 0 252522 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 254122 0 254178 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 255686 0 255742 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 257342 0 257398 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 142066 0 142122 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 151634 0 151690 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 153290 0 153346 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 154854 0 154910 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 164514 0 164570 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 175646 0 175702 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 178866 0 178922 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 180430 0 180486 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 182086 0 182142 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 183650 0 183706 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 185306 0 185362 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 186870 0 186926 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 190090 0 190146 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 191654 0 191710 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 193310 0 193366 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 196438 0 196494 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 198094 0 198150 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 201314 0 201370 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 202878 0 202934 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 204442 0 204498 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 206098 0 206154 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 207662 0 207718 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 212446 0 212502 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 215666 0 215722 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 217782 0 217838 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 221002 0 221058 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 224222 0 224278 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 225786 0 225842 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 229006 0 229062 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 230662 0 230718 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 232226 0 232282 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 238666 0 238722 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 243450 0 243506 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 249798 0 249854 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 251454 0 251510 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 253018 0 253074 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 254674 0 254730 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 257802 0 257858 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 259458 0 259514 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 261022 0 261078 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 196990 0 197046 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 200210 0 200266 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 201774 0 201830 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 203430 0 203486 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 206650 0 206706 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 214654 0 214710 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 216218 0 216274 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 249968 2128 250288 262256 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 262256 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 262256 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 262256 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 262256 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 262256 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 262256 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 262256 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 262256 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 234608 2128 234928 262256 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 262256 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 262256 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 262256 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 262256 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 262256 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 262256 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 262256 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 250628 2176 250948 262208 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 262208 6 vccd2
port 626 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 262208 6 vccd2
port 627 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 262208 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 262208 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 262208 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 262208 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 262208 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 262208 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 235268 2176 235588 262208 6 vssd2
port 634 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 262208 6 vssd2
port 635 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 262208 6 vssd2
port 636 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 262208 6 vssd2
port 637 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 262208 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 262208 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 262208 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 262208 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 251288 2176 251608 262208 6 vdda1
port 642 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 262208 6 vdda1
port 643 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 262208 6 vdda1
port 644 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 262208 6 vdda1
port 645 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 262208 6 vdda1
port 646 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 262208 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 262208 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 262208 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 262208 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 235928 2176 236248 262208 6 vssa1
port 651 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 262208 6 vssa1
port 652 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 262208 6 vssa1
port 653 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 262208 6 vssa1
port 654 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 262208 6 vssa1
port 655 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 262208 6 vssa1
port 656 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 262208 6 vssa1
port 657 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 262208 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 251948 2176 252268 262208 6 vdda2
port 659 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 262208 6 vdda2
port 660 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 262208 6 vdda2
port 661 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 262208 6 vdda2
port 662 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 262208 6 vdda2
port 663 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 262208 6 vdda2
port 664 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 262208 6 vdda2
port 665 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 262208 6 vdda2
port 666 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 262208 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 236588 2176 236908 262208 6 vssa2
port 668 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 262208 6 vssa2
port 669 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 262208 6 vssa2
port 670 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 262208 6 vssa2
port 671 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 262208 6 vssa2
port 672 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 262208 6 vssa2
port 673 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 262208 6 vssa2
port 674 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 262208 6 vssa2
port 675 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 262521 264665
string LEFview TRUE
string GDS_FILE /project/openlane/axi_dma/runs/axi_dma/results/magic/axi_dma.gds
string GDS_END 98131030
string GDS_START 1183208
<< end >>

