magic
tech sky130A
magscale 1 2
timestamp 1622715337
<< obsli1 >>
rect 1104 2159 179584 180625
<< obsm1 >>
rect 198 1980 180582 180656
<< metal2 >>
rect 754 182088 810 182888
rect 2318 182088 2374 182888
rect 3882 182088 3938 182888
rect 5446 182088 5502 182888
rect 7010 182088 7066 182888
rect 8666 182088 8722 182888
rect 10230 182088 10286 182888
rect 11794 182088 11850 182888
rect 13358 182088 13414 182888
rect 15014 182088 15070 182888
rect 16578 182088 16634 182888
rect 18142 182088 18198 182888
rect 19706 182088 19762 182888
rect 21362 182088 21418 182888
rect 22926 182088 22982 182888
rect 24490 182088 24546 182888
rect 26054 182088 26110 182888
rect 27710 182088 27766 182888
rect 29274 182088 29330 182888
rect 30838 182088 30894 182888
rect 32402 182088 32458 182888
rect 33966 182088 34022 182888
rect 35622 182088 35678 182888
rect 37186 182088 37242 182888
rect 38750 182088 38806 182888
rect 40314 182088 40370 182888
rect 41970 182088 42026 182888
rect 43534 182088 43590 182888
rect 45098 182088 45154 182888
rect 46662 182088 46718 182888
rect 48318 182088 48374 182888
rect 49882 182088 49938 182888
rect 51446 182088 51502 182888
rect 53010 182088 53066 182888
rect 54666 182088 54722 182888
rect 56230 182088 56286 182888
rect 57794 182088 57850 182888
rect 59358 182088 59414 182888
rect 61014 182088 61070 182888
rect 62578 182088 62634 182888
rect 64142 182088 64198 182888
rect 65706 182088 65762 182888
rect 67270 182088 67326 182888
rect 68926 182088 68982 182888
rect 70490 182088 70546 182888
rect 72054 182088 72110 182888
rect 73618 182088 73674 182888
rect 75274 182088 75330 182888
rect 76838 182088 76894 182888
rect 78402 182088 78458 182888
rect 79966 182088 80022 182888
rect 81622 182088 81678 182888
rect 83186 182088 83242 182888
rect 84750 182088 84806 182888
rect 86314 182088 86370 182888
rect 87970 182088 88026 182888
rect 89534 182088 89590 182888
rect 91098 182088 91154 182888
rect 92662 182088 92718 182888
rect 94226 182088 94282 182888
rect 95882 182088 95938 182888
rect 97446 182088 97502 182888
rect 99010 182088 99066 182888
rect 100574 182088 100630 182888
rect 102230 182088 102286 182888
rect 103794 182088 103850 182888
rect 105358 182088 105414 182888
rect 106922 182088 106978 182888
rect 108578 182088 108634 182888
rect 110142 182088 110198 182888
rect 111706 182088 111762 182888
rect 113270 182088 113326 182888
rect 114926 182088 114982 182888
rect 116490 182088 116546 182888
rect 118054 182088 118110 182888
rect 119618 182088 119674 182888
rect 121274 182088 121330 182888
rect 122838 182088 122894 182888
rect 124402 182088 124458 182888
rect 125966 182088 126022 182888
rect 127530 182088 127586 182888
rect 129186 182088 129242 182888
rect 130750 182088 130806 182888
rect 132314 182088 132370 182888
rect 133878 182088 133934 182888
rect 135534 182088 135590 182888
rect 137098 182088 137154 182888
rect 138662 182088 138718 182888
rect 140226 182088 140282 182888
rect 141882 182088 141938 182888
rect 143446 182088 143502 182888
rect 145010 182088 145066 182888
rect 146574 182088 146630 182888
rect 148230 182088 148286 182888
rect 149794 182088 149850 182888
rect 151358 182088 151414 182888
rect 152922 182088 152978 182888
rect 154486 182088 154542 182888
rect 156142 182088 156198 182888
rect 157706 182088 157762 182888
rect 159270 182088 159326 182888
rect 160834 182088 160890 182888
rect 162490 182088 162546 182888
rect 164054 182088 164110 182888
rect 165618 182088 165674 182888
rect 167182 182088 167238 182888
rect 168838 182088 168894 182888
rect 170402 182088 170458 182888
rect 171966 182088 172022 182888
rect 173530 182088 173586 182888
rect 175186 182088 175242 182888
rect 176750 182088 176806 182888
rect 178314 182088 178370 182888
rect 179878 182088 179934 182888
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43350 0 43406 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45926 0 45982 800
rect 46294 0 46350 800
rect 46662 0 46718 800
rect 47030 0 47086 800
rect 47398 0 47454 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48502 0 48558 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51814 0 51870 800
rect 52182 0 52238 800
rect 52550 0 52606 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54390 0 54446 800
rect 54758 0 54814 800
rect 55126 0 55182 800
rect 55494 0 55550 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57702 0 57758 800
rect 58070 0 58126 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59174 0 59230 800
rect 59542 0 59598 800
rect 59910 0 59966 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70582 0 70638 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72514 0 72570 800
rect 72882 0 72938 800
rect 73250 0 73306 800
rect 73618 0 73674 800
rect 73986 0 74042 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 75090 0 75146 800
rect 75458 0 75514 800
rect 75826 0 75882 800
rect 76194 0 76250 800
rect 76562 0 76618 800
rect 76930 0 76986 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 78034 0 78090 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79138 0 79194 800
rect 79506 0 79562 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80610 0 80666 800
rect 80978 0 81034 800
rect 81346 0 81402 800
rect 81714 0 81770 800
rect 82082 0 82138 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83186 0 83242 800
rect 83554 0 83610 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87234 0 87290 800
rect 87602 0 87658 800
rect 87970 0 88026 800
rect 88338 0 88394 800
rect 88706 0 88762 800
rect 89074 0 89130 800
rect 89442 0 89498 800
rect 89810 0 89866 800
rect 90178 0 90234 800
rect 90546 0 90602 800
rect 90914 0 90970 800
rect 91282 0 91338 800
rect 91650 0 91706 800
rect 92018 0 92074 800
rect 92386 0 92442 800
rect 92754 0 92810 800
rect 93122 0 93178 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94962 0 95018 800
rect 95330 0 95386 800
rect 95698 0 95754 800
rect 96066 0 96122 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97170 0 97226 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100114 0 100170 800
rect 100482 0 100538 800
rect 100850 0 100906 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102690 0 102746 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108210 0 108266 800
rect 108670 0 108726 800
rect 109038 0 109094 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110142 0 110198 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 113086 0 113142 800
rect 113454 0 113510 800
rect 113822 0 113878 800
rect 114190 0 114246 800
rect 114558 0 114614 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116766 0 116822 800
rect 117134 0 117190 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118238 0 118294 800
rect 118606 0 118662 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124494 0 124550 800
rect 124862 0 124918 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126702 0 126758 800
rect 127070 0 127126 800
rect 127438 0 127494 800
rect 127806 0 127862 800
rect 128174 0 128230 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129278 0 129334 800
rect 129646 0 129702 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131118 0 131174 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132222 0 132278 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133694 0 133750 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134798 0 134854 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137374 0 137430 800
rect 137742 0 137798 800
rect 138110 0 138166 800
rect 138478 0 138534 800
rect 138846 0 138902 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140318 0 140374 800
rect 140686 0 140742 800
rect 141054 0 141110 800
rect 141422 0 141478 800
rect 141790 0 141846 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 143998 0 144054 800
rect 144366 0 144422 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
rect 180154 0 180210 800
rect 180522 0 180578 800
<< obsm2 >>
rect 204 182032 698 182088
rect 866 182032 2262 182088
rect 2430 182032 3826 182088
rect 3994 182032 5390 182088
rect 5558 182032 6954 182088
rect 7122 182032 8610 182088
rect 8778 182032 10174 182088
rect 10342 182032 11738 182088
rect 11906 182032 13302 182088
rect 13470 182032 14958 182088
rect 15126 182032 16522 182088
rect 16690 182032 18086 182088
rect 18254 182032 19650 182088
rect 19818 182032 21306 182088
rect 21474 182032 22870 182088
rect 23038 182032 24434 182088
rect 24602 182032 25998 182088
rect 26166 182032 27654 182088
rect 27822 182032 29218 182088
rect 29386 182032 30782 182088
rect 30950 182032 32346 182088
rect 32514 182032 33910 182088
rect 34078 182032 35566 182088
rect 35734 182032 37130 182088
rect 37298 182032 38694 182088
rect 38862 182032 40258 182088
rect 40426 182032 41914 182088
rect 42082 182032 43478 182088
rect 43646 182032 45042 182088
rect 45210 182032 46606 182088
rect 46774 182032 48262 182088
rect 48430 182032 49826 182088
rect 49994 182032 51390 182088
rect 51558 182032 52954 182088
rect 53122 182032 54610 182088
rect 54778 182032 56174 182088
rect 56342 182032 57738 182088
rect 57906 182032 59302 182088
rect 59470 182032 60958 182088
rect 61126 182032 62522 182088
rect 62690 182032 64086 182088
rect 64254 182032 65650 182088
rect 65818 182032 67214 182088
rect 67382 182032 68870 182088
rect 69038 182032 70434 182088
rect 70602 182032 71998 182088
rect 72166 182032 73562 182088
rect 73730 182032 75218 182088
rect 75386 182032 76782 182088
rect 76950 182032 78346 182088
rect 78514 182032 79910 182088
rect 80078 182032 81566 182088
rect 81734 182032 83130 182088
rect 83298 182032 84694 182088
rect 84862 182032 86258 182088
rect 86426 182032 87914 182088
rect 88082 182032 89478 182088
rect 89646 182032 91042 182088
rect 91210 182032 92606 182088
rect 92774 182032 94170 182088
rect 94338 182032 95826 182088
rect 95994 182032 97390 182088
rect 97558 182032 98954 182088
rect 99122 182032 100518 182088
rect 100686 182032 102174 182088
rect 102342 182032 103738 182088
rect 103906 182032 105302 182088
rect 105470 182032 106866 182088
rect 107034 182032 108522 182088
rect 108690 182032 110086 182088
rect 110254 182032 111650 182088
rect 111818 182032 113214 182088
rect 113382 182032 114870 182088
rect 115038 182032 116434 182088
rect 116602 182032 117998 182088
rect 118166 182032 119562 182088
rect 119730 182032 121218 182088
rect 121386 182032 122782 182088
rect 122950 182032 124346 182088
rect 124514 182032 125910 182088
rect 126078 182032 127474 182088
rect 127642 182032 129130 182088
rect 129298 182032 130694 182088
rect 130862 182032 132258 182088
rect 132426 182032 133822 182088
rect 133990 182032 135478 182088
rect 135646 182032 137042 182088
rect 137210 182032 138606 182088
rect 138774 182032 140170 182088
rect 140338 182032 141826 182088
rect 141994 182032 143390 182088
rect 143558 182032 144954 182088
rect 145122 182032 146518 182088
rect 146686 182032 148174 182088
rect 148342 182032 149738 182088
rect 149906 182032 151302 182088
rect 151470 182032 152866 182088
rect 153034 182032 154430 182088
rect 154598 182032 156086 182088
rect 156254 182032 157650 182088
rect 157818 182032 159214 182088
rect 159382 182032 160778 182088
rect 160946 182032 162434 182088
rect 162602 182032 163998 182088
rect 164166 182032 165562 182088
rect 165730 182032 167126 182088
rect 167294 182032 168782 182088
rect 168950 182032 170346 182088
rect 170514 182032 171910 182088
rect 172078 182032 173474 182088
rect 173642 182032 175130 182088
rect 175298 182032 176694 182088
rect 176862 182032 178258 182088
rect 178426 182032 179822 182088
rect 179990 182032 180576 182088
rect 204 856 180576 182032
rect 314 800 514 856
rect 682 800 882 856
rect 1050 800 1250 856
rect 1418 800 1618 856
rect 1786 800 1986 856
rect 2154 800 2354 856
rect 2522 800 2722 856
rect 2890 800 3090 856
rect 3258 800 3458 856
rect 3626 800 3826 856
rect 3994 800 4194 856
rect 4362 800 4562 856
rect 4730 800 4930 856
rect 5098 800 5298 856
rect 5466 800 5666 856
rect 5834 800 6034 856
rect 6202 800 6402 856
rect 6570 800 6770 856
rect 6938 800 7138 856
rect 7306 800 7506 856
rect 7674 800 7874 856
rect 8042 800 8242 856
rect 8410 800 8610 856
rect 8778 800 8978 856
rect 9146 800 9346 856
rect 9514 800 9714 856
rect 9882 800 10082 856
rect 10250 800 10450 856
rect 10618 800 10818 856
rect 10986 800 11186 856
rect 11354 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12658 856
rect 12826 800 13026 856
rect 13194 800 13394 856
rect 13562 800 13762 856
rect 13930 800 14130 856
rect 14298 800 14498 856
rect 14666 800 14866 856
rect 15034 800 15234 856
rect 15402 800 15602 856
rect 15770 800 15970 856
rect 16138 800 16338 856
rect 16506 800 16706 856
rect 16874 800 17074 856
rect 17242 800 17442 856
rect 17610 800 17810 856
rect 17978 800 18178 856
rect 18346 800 18546 856
rect 18714 800 18914 856
rect 19082 800 19282 856
rect 19450 800 19650 856
rect 19818 800 20018 856
rect 20186 800 20386 856
rect 20554 800 20754 856
rect 20922 800 21122 856
rect 21290 800 21490 856
rect 21658 800 21858 856
rect 22026 800 22226 856
rect 22394 800 22594 856
rect 22762 800 22962 856
rect 23130 800 23330 856
rect 23498 800 23698 856
rect 23866 800 24066 856
rect 24234 800 24434 856
rect 24602 800 24802 856
rect 24970 800 25170 856
rect 25338 800 25538 856
rect 25706 800 25906 856
rect 26074 800 26274 856
rect 26442 800 26642 856
rect 26810 800 27010 856
rect 27178 800 27378 856
rect 27546 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28482 856
rect 28650 800 28850 856
rect 29018 800 29218 856
rect 29386 800 29586 856
rect 29754 800 29954 856
rect 30122 800 30322 856
rect 30490 800 30690 856
rect 30858 800 31058 856
rect 31226 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32530 856
rect 32698 800 32898 856
rect 33066 800 33266 856
rect 33434 800 33634 856
rect 33802 800 34002 856
rect 34170 800 34370 856
rect 34538 800 34738 856
rect 34906 800 35106 856
rect 35274 800 35474 856
rect 35642 800 35842 856
rect 36010 800 36302 856
rect 36470 800 36670 856
rect 36838 800 37038 856
rect 37206 800 37406 856
rect 37574 800 37774 856
rect 37942 800 38142 856
rect 38310 800 38510 856
rect 38678 800 38878 856
rect 39046 800 39246 856
rect 39414 800 39614 856
rect 39782 800 39982 856
rect 40150 800 40350 856
rect 40518 800 40718 856
rect 40886 800 41086 856
rect 41254 800 41454 856
rect 41622 800 41822 856
rect 41990 800 42190 856
rect 42358 800 42558 856
rect 42726 800 42926 856
rect 43094 800 43294 856
rect 43462 800 43662 856
rect 43830 800 44030 856
rect 44198 800 44398 856
rect 44566 800 44766 856
rect 44934 800 45134 856
rect 45302 800 45502 856
rect 45670 800 45870 856
rect 46038 800 46238 856
rect 46406 800 46606 856
rect 46774 800 46974 856
rect 47142 800 47342 856
rect 47510 800 47710 856
rect 47878 800 48078 856
rect 48246 800 48446 856
rect 48614 800 48814 856
rect 48982 800 49182 856
rect 49350 800 49550 856
rect 49718 800 49918 856
rect 50086 800 50286 856
rect 50454 800 50654 856
rect 50822 800 51022 856
rect 51190 800 51390 856
rect 51558 800 51758 856
rect 51926 800 52126 856
rect 52294 800 52494 856
rect 52662 800 52862 856
rect 53030 800 53230 856
rect 53398 800 53598 856
rect 53766 800 53966 856
rect 54134 800 54334 856
rect 54502 800 54702 856
rect 54870 800 55070 856
rect 55238 800 55438 856
rect 55606 800 55806 856
rect 55974 800 56174 856
rect 56342 800 56542 856
rect 56710 800 56910 856
rect 57078 800 57278 856
rect 57446 800 57646 856
rect 57814 800 58014 856
rect 58182 800 58382 856
rect 58550 800 58750 856
rect 58918 800 59118 856
rect 59286 800 59486 856
rect 59654 800 59854 856
rect 60022 800 60222 856
rect 60390 800 60590 856
rect 60758 800 60958 856
rect 61126 800 61326 856
rect 61494 800 61694 856
rect 61862 800 62062 856
rect 62230 800 62430 856
rect 62598 800 62798 856
rect 62966 800 63166 856
rect 63334 800 63534 856
rect 63702 800 63902 856
rect 64070 800 64270 856
rect 64438 800 64638 856
rect 64806 800 65006 856
rect 65174 800 65374 856
rect 65542 800 65742 856
rect 65910 800 66110 856
rect 66278 800 66478 856
rect 66646 800 66846 856
rect 67014 800 67214 856
rect 67382 800 67582 856
rect 67750 800 67950 856
rect 68118 800 68318 856
rect 68486 800 68686 856
rect 68854 800 69054 856
rect 69222 800 69422 856
rect 69590 800 69790 856
rect 69958 800 70158 856
rect 70326 800 70526 856
rect 70694 800 70894 856
rect 71062 800 71262 856
rect 71430 800 71630 856
rect 71798 800 71998 856
rect 72166 800 72458 856
rect 72626 800 72826 856
rect 72994 800 73194 856
rect 73362 800 73562 856
rect 73730 800 73930 856
rect 74098 800 74298 856
rect 74466 800 74666 856
rect 74834 800 75034 856
rect 75202 800 75402 856
rect 75570 800 75770 856
rect 75938 800 76138 856
rect 76306 800 76506 856
rect 76674 800 76874 856
rect 77042 800 77242 856
rect 77410 800 77610 856
rect 77778 800 77978 856
rect 78146 800 78346 856
rect 78514 800 78714 856
rect 78882 800 79082 856
rect 79250 800 79450 856
rect 79618 800 79818 856
rect 79986 800 80186 856
rect 80354 800 80554 856
rect 80722 800 80922 856
rect 81090 800 81290 856
rect 81458 800 81658 856
rect 81826 800 82026 856
rect 82194 800 82394 856
rect 82562 800 82762 856
rect 82930 800 83130 856
rect 83298 800 83498 856
rect 83666 800 83866 856
rect 84034 800 84234 856
rect 84402 800 84602 856
rect 84770 800 84970 856
rect 85138 800 85338 856
rect 85506 800 85706 856
rect 85874 800 86074 856
rect 86242 800 86442 856
rect 86610 800 86810 856
rect 86978 800 87178 856
rect 87346 800 87546 856
rect 87714 800 87914 856
rect 88082 800 88282 856
rect 88450 800 88650 856
rect 88818 800 89018 856
rect 89186 800 89386 856
rect 89554 800 89754 856
rect 89922 800 90122 856
rect 90290 800 90490 856
rect 90658 800 90858 856
rect 91026 800 91226 856
rect 91394 800 91594 856
rect 91762 800 91962 856
rect 92130 800 92330 856
rect 92498 800 92698 856
rect 92866 800 93066 856
rect 93234 800 93434 856
rect 93602 800 93802 856
rect 93970 800 94170 856
rect 94338 800 94538 856
rect 94706 800 94906 856
rect 95074 800 95274 856
rect 95442 800 95642 856
rect 95810 800 96010 856
rect 96178 800 96378 856
rect 96546 800 96746 856
rect 96914 800 97114 856
rect 97282 800 97482 856
rect 97650 800 97850 856
rect 98018 800 98218 856
rect 98386 800 98586 856
rect 98754 800 98954 856
rect 99122 800 99322 856
rect 99490 800 99690 856
rect 99858 800 100058 856
rect 100226 800 100426 856
rect 100594 800 100794 856
rect 100962 800 101162 856
rect 101330 800 101530 856
rect 101698 800 101898 856
rect 102066 800 102266 856
rect 102434 800 102634 856
rect 102802 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104474 856
rect 104642 800 104842 856
rect 105010 800 105210 856
rect 105378 800 105578 856
rect 105746 800 105946 856
rect 106114 800 106314 856
rect 106482 800 106682 856
rect 106850 800 107050 856
rect 107218 800 107418 856
rect 107586 800 107786 856
rect 107954 800 108154 856
rect 108322 800 108614 856
rect 108782 800 108982 856
rect 109150 800 109350 856
rect 109518 800 109718 856
rect 109886 800 110086 856
rect 110254 800 110454 856
rect 110622 800 110822 856
rect 110990 800 111190 856
rect 111358 800 111558 856
rect 111726 800 111926 856
rect 112094 800 112294 856
rect 112462 800 112662 856
rect 112830 800 113030 856
rect 113198 800 113398 856
rect 113566 800 113766 856
rect 113934 800 114134 856
rect 114302 800 114502 856
rect 114670 800 114870 856
rect 115038 800 115238 856
rect 115406 800 115606 856
rect 115774 800 115974 856
rect 116142 800 116342 856
rect 116510 800 116710 856
rect 116878 800 117078 856
rect 117246 800 117446 856
rect 117614 800 117814 856
rect 117982 800 118182 856
rect 118350 800 118550 856
rect 118718 800 118918 856
rect 119086 800 119286 856
rect 119454 800 119654 856
rect 119822 800 120022 856
rect 120190 800 120390 856
rect 120558 800 120758 856
rect 120926 800 121126 856
rect 121294 800 121494 856
rect 121662 800 121862 856
rect 122030 800 122230 856
rect 122398 800 122598 856
rect 122766 800 122966 856
rect 123134 800 123334 856
rect 123502 800 123702 856
rect 123870 800 124070 856
rect 124238 800 124438 856
rect 124606 800 124806 856
rect 124974 800 125174 856
rect 125342 800 125542 856
rect 125710 800 125910 856
rect 126078 800 126278 856
rect 126446 800 126646 856
rect 126814 800 127014 856
rect 127182 800 127382 856
rect 127550 800 127750 856
rect 127918 800 128118 856
rect 128286 800 128486 856
rect 128654 800 128854 856
rect 129022 800 129222 856
rect 129390 800 129590 856
rect 129758 800 129958 856
rect 130126 800 130326 856
rect 130494 800 130694 856
rect 130862 800 131062 856
rect 131230 800 131430 856
rect 131598 800 131798 856
rect 131966 800 132166 856
rect 132334 800 132534 856
rect 132702 800 132902 856
rect 133070 800 133270 856
rect 133438 800 133638 856
rect 133806 800 134006 856
rect 134174 800 134374 856
rect 134542 800 134742 856
rect 134910 800 135110 856
rect 135278 800 135478 856
rect 135646 800 135846 856
rect 136014 800 136214 856
rect 136382 800 136582 856
rect 136750 800 136950 856
rect 137118 800 137318 856
rect 137486 800 137686 856
rect 137854 800 138054 856
rect 138222 800 138422 856
rect 138590 800 138790 856
rect 138958 800 139158 856
rect 139326 800 139526 856
rect 139694 800 139894 856
rect 140062 800 140262 856
rect 140430 800 140630 856
rect 140798 800 140998 856
rect 141166 800 141366 856
rect 141534 800 141734 856
rect 141902 800 142102 856
rect 142270 800 142470 856
rect 142638 800 142838 856
rect 143006 800 143206 856
rect 143374 800 143574 856
rect 143742 800 143942 856
rect 144110 800 144310 856
rect 144478 800 144770 856
rect 144938 800 145138 856
rect 145306 800 145506 856
rect 145674 800 145874 856
rect 146042 800 146242 856
rect 146410 800 146610 856
rect 146778 800 146978 856
rect 147146 800 147346 856
rect 147514 800 147714 856
rect 147882 800 148082 856
rect 148250 800 148450 856
rect 148618 800 148818 856
rect 148986 800 149186 856
rect 149354 800 149554 856
rect 149722 800 149922 856
rect 150090 800 150290 856
rect 150458 800 150658 856
rect 150826 800 151026 856
rect 151194 800 151394 856
rect 151562 800 151762 856
rect 151930 800 152130 856
rect 152298 800 152498 856
rect 152666 800 152866 856
rect 153034 800 153234 856
rect 153402 800 153602 856
rect 153770 800 153970 856
rect 154138 800 154338 856
rect 154506 800 154706 856
rect 154874 800 155074 856
rect 155242 800 155442 856
rect 155610 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156546 856
rect 156714 800 156914 856
rect 157082 800 157282 856
rect 157450 800 157650 856
rect 157818 800 158018 856
rect 158186 800 158386 856
rect 158554 800 158754 856
rect 158922 800 159122 856
rect 159290 800 159490 856
rect 159658 800 159858 856
rect 160026 800 160226 856
rect 160394 800 160594 856
rect 160762 800 160962 856
rect 161130 800 161330 856
rect 161498 800 161698 856
rect 161866 800 162066 856
rect 162234 800 162434 856
rect 162602 800 162802 856
rect 162970 800 163170 856
rect 163338 800 163538 856
rect 163706 800 163906 856
rect 164074 800 164274 856
rect 164442 800 164642 856
rect 164810 800 165010 856
rect 165178 800 165378 856
rect 165546 800 165746 856
rect 165914 800 166114 856
rect 166282 800 166482 856
rect 166650 800 166850 856
rect 167018 800 167218 856
rect 167386 800 167586 856
rect 167754 800 167954 856
rect 168122 800 168322 856
rect 168490 800 168690 856
rect 168858 800 169058 856
rect 169226 800 169426 856
rect 169594 800 169794 856
rect 169962 800 170162 856
rect 170330 800 170530 856
rect 170698 800 170898 856
rect 171066 800 171266 856
rect 171434 800 171634 856
rect 171802 800 172002 856
rect 172170 800 172370 856
rect 172538 800 172738 856
rect 172906 800 173106 856
rect 173274 800 173474 856
rect 173642 800 173842 856
rect 174010 800 174210 856
rect 174378 800 174578 856
rect 174746 800 174946 856
rect 175114 800 175314 856
rect 175482 800 175682 856
rect 175850 800 176050 856
rect 176218 800 176418 856
rect 176586 800 176786 856
rect 176954 800 177154 856
rect 177322 800 177522 856
rect 177690 800 177890 856
rect 178058 800 178258 856
rect 178426 800 178626 856
rect 178794 800 178994 856
rect 179162 800 179362 856
rect 179530 800 179730 856
rect 179898 800 180098 856
rect 180266 800 180466 856
<< metal3 >>
rect 0 137096 800 137216
rect 179944 91400 180744 91520
rect 0 45704 800 45824
<< obsm3 >>
rect 800 137296 179944 180641
rect 880 137016 179944 137296
rect 800 91600 179944 137016
rect 800 91320 179864 91600
rect 800 45904 179944 91320
rect 880 45624 179944 45904
rect 800 2143 179944 45624
<< metal4 >>
rect 4208 2128 4528 180656
rect 4868 2176 5188 180608
rect 5528 2176 5848 180608
rect 6188 2176 6508 180608
rect 19568 2128 19888 180656
rect 20228 2176 20548 180608
rect 20888 2176 21208 180608
rect 21548 2176 21868 180608
rect 34928 2128 35248 180656
rect 35588 2176 35908 180608
rect 36248 2176 36568 180608
rect 36908 2176 37228 180608
rect 50288 2128 50608 180656
rect 50948 2176 51268 180608
rect 51608 2176 51928 180608
rect 52268 2176 52588 180608
rect 65648 2128 65968 180656
rect 66308 2176 66628 180608
rect 66968 2176 67288 180608
rect 67628 2176 67948 180608
rect 81008 2128 81328 180656
rect 81668 2176 81988 180608
rect 82328 2176 82648 180608
rect 82988 2176 83308 180608
rect 96368 2128 96688 180656
rect 97028 2176 97348 180608
rect 97688 2176 98008 180608
rect 98348 2176 98668 180608
rect 111728 2128 112048 180656
rect 112388 2176 112708 180608
rect 113048 2176 113368 180608
rect 113708 2176 114028 180608
rect 127088 2128 127408 180656
rect 127748 2176 128068 180608
rect 128408 2176 128728 180608
rect 129068 2176 129388 180608
rect 142448 2128 142768 180656
rect 143108 2176 143428 180608
rect 143768 2176 144088 180608
rect 144428 2176 144748 180608
rect 157808 2128 158128 180656
rect 158468 2176 158788 180608
rect 159128 2176 159448 180608
rect 159788 2176 160108 180608
rect 173168 2128 173488 180656
rect 173828 2176 174148 180608
rect 174488 2176 174808 180608
rect 175148 2176 175468 180608
<< obsm4 >>
rect 19379 2483 19488 146437
rect 19968 2483 20148 146437
rect 20628 2483 20808 146437
rect 21288 2483 21468 146437
rect 21948 2483 34848 146437
rect 35328 2483 35508 146437
rect 35988 2483 36168 146437
rect 36648 2483 36828 146437
rect 37308 2483 50208 146437
rect 50688 2483 50868 146437
rect 51348 2483 51528 146437
rect 52008 2483 52188 146437
rect 52668 2483 65568 146437
rect 66048 2483 66228 146437
rect 66708 2483 66888 146437
rect 67368 2483 67548 146437
rect 68028 2483 80928 146437
rect 81408 2483 81588 146437
rect 82068 2483 82248 146437
rect 82728 2483 82908 146437
rect 83388 2483 96288 146437
rect 96768 2483 96948 146437
rect 97428 2483 97608 146437
rect 98088 2483 98268 146437
rect 98748 2483 111648 146437
rect 112128 2483 112308 146437
rect 112788 2483 112968 146437
rect 113448 2483 113628 146437
rect 114108 2483 125429 146437
<< labels >>
rlabel metal2 s 754 182088 810 182888 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 48318 182088 48374 182888 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 53010 182088 53066 182888 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57794 182088 57850 182888 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 62578 182088 62634 182888 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 67270 182088 67326 182888 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 72054 182088 72110 182888 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 76838 182088 76894 182888 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 81622 182088 81678 182888 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 86314 182088 86370 182888 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 91098 182088 91154 182888 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5446 182088 5502 182888 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 95882 182088 95938 182888 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 100574 182088 100630 182888 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 105358 182088 105414 182888 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 110142 182088 110198 182888 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 114926 182088 114982 182888 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 119618 182088 119674 182888 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 124402 182088 124458 182888 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 129186 182088 129242 182888 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 133878 182088 133934 182888 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 138662 182088 138718 182888 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10230 182088 10286 182888 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 143446 182088 143502 182888 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 148230 182088 148286 182888 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 152922 182088 152978 182888 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 157706 182088 157762 182888 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 162490 182088 162546 182888 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 167182 182088 167238 182888 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 171966 182088 172022 182888 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 176750 182088 176806 182888 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 15014 182088 15070 182888 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 19706 182088 19762 182888 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 24490 182088 24546 182888 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 29274 182088 29330 182888 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 33966 182088 34022 182888 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 38750 182088 38806 182888 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 43534 182088 43590 182888 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2318 182088 2374 182888 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 49882 182088 49938 182888 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 54666 182088 54722 182888 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 59358 182088 59414 182888 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 64142 182088 64198 182888 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68926 182088 68982 182888 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 73618 182088 73674 182888 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 78402 182088 78458 182888 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 83186 182088 83242 182888 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 87970 182088 88026 182888 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 92662 182088 92718 182888 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7010 182088 7066 182888 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 97446 182088 97502 182888 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 102230 182088 102286 182888 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 106922 182088 106978 182888 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 111706 182088 111762 182888 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 116490 182088 116546 182888 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 121274 182088 121330 182888 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 125966 182088 126022 182888 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 130750 182088 130806 182888 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 135534 182088 135590 182888 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 140226 182088 140282 182888 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11794 182088 11850 182888 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 145010 182088 145066 182888 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 149794 182088 149850 182888 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 154486 182088 154542 182888 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 159270 182088 159326 182888 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 164054 182088 164110 182888 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 168838 182088 168894 182888 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 173530 182088 173586 182888 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 178314 182088 178370 182888 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 16578 182088 16634 182888 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21362 182088 21418 182888 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 26054 182088 26110 182888 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 30838 182088 30894 182888 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35622 182088 35678 182888 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 40314 182088 40370 182888 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 45098 182088 45154 182888 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3882 182088 3938 182888 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 51446 182088 51502 182888 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 56230 182088 56286 182888 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 61014 182088 61070 182888 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 65706 182088 65762 182888 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 70490 182088 70546 182888 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 75274 182088 75330 182888 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 79966 182088 80022 182888 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 84750 182088 84806 182888 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 89534 182088 89590 182888 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 94226 182088 94282 182888 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8666 182088 8722 182888 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 99010 182088 99066 182888 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 103794 182088 103850 182888 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 108578 182088 108634 182888 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 113270 182088 113326 182888 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 118054 182088 118110 182888 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 122838 182088 122894 182888 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 127530 182088 127586 182888 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 132314 182088 132370 182888 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 137098 182088 137154 182888 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 141882 182088 141938 182888 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13358 182088 13414 182888 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 146574 182088 146630 182888 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 151358 182088 151414 182888 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 156142 182088 156198 182888 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 160834 182088 160890 182888 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 165618 182088 165674 182888 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 170402 182088 170458 182888 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 175186 182088 175242 182888 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 179878 182088 179934 182888 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 18142 182088 18198 182888 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 22926 182088 22982 182888 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 27710 182088 27766 182888 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32402 182088 32458 182888 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37186 182088 37242 182888 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 41970 182088 42026 182888 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46662 182088 46718 182888 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 179944 91400 180744 91520 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 0 137096 800 137216 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 150346 0 150402 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 151450 0 151506 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 169114 0 169170 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 174634 0 174690 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 180154 0 180210 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 121550 0 121606 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 138110 0 138166 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 141422 0 141478 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 142526 0 142582 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 149242 0 149298 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 2410 0 2466 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 157808 2128 158128 180656 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 180656 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 180656 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 180656 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 180656 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 180656 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 180656 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 180656 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 180656 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 180656 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 180656 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 180656 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 180608 6 vccd2
port 620 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 180608 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 180608 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 180608 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 180608 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 180608 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 180608 6 vssd2
port 626 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 180608 6 vssd2
port 627 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 180608 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 180608 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 180608 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 180608 6 vssd2
port 631 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 180608 6 vdda1
port 632 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 180608 6 vdda1
port 633 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 180608 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 180608 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 180608 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 180608 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 180608 6 vssa1
port 638 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 180608 6 vssa1
port 639 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 180608 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 180608 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 180608 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 180608 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 180608 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 180608 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 180608 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 180608 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 180608 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 180608 6 vdda2
port 649 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 180608 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 180608 6 vssa2
port 651 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 180608 6 vssa2
port 652 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 180608 6 vssa2
port 653 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 180608 6 vssa2
port 654 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 180608 6 vssa2
port 655 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180744 182888
string LEFview TRUE
string GDS_FILE /project/openlane/axi_dma/runs/axi_dma/results/magic/axi_dma.gds
string GDS_END 56515138
string GDS_START 1195668
<< end >>

