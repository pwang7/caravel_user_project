magic
tech sky130A
magscale 1 2
timestamp 1623901464
<< obsli1 >>
rect 1104 1377 260084 261137
<< obsm1 >>
rect 198 1096 260898 261168
<< metal2 >>
rect 1122 262535 1178 263335
rect 3330 262535 3386 263335
rect 5630 262535 5686 263335
rect 7930 262535 7986 263335
rect 10138 262535 10194 263335
rect 12438 262535 12494 263335
rect 14738 262535 14794 263335
rect 16946 262535 17002 263335
rect 19246 262535 19302 263335
rect 21546 262535 21602 263335
rect 23754 262535 23810 263335
rect 26054 262535 26110 263335
rect 28354 262535 28410 263335
rect 30562 262535 30618 263335
rect 32862 262535 32918 263335
rect 35162 262535 35218 263335
rect 37370 262535 37426 263335
rect 39670 262535 39726 263335
rect 41970 262535 42026 263335
rect 44270 262535 44326 263335
rect 46478 262535 46534 263335
rect 48778 262535 48834 263335
rect 51078 262535 51134 263335
rect 53286 262535 53342 263335
rect 55586 262535 55642 263335
rect 57886 262535 57942 263335
rect 60094 262535 60150 263335
rect 62394 262535 62450 263335
rect 64694 262535 64750 263335
rect 66902 262535 66958 263335
rect 69202 262535 69258 263335
rect 71502 262535 71558 263335
rect 73710 262535 73766 263335
rect 76010 262535 76066 263335
rect 78310 262535 78366 263335
rect 80610 262535 80666 263335
rect 82818 262535 82874 263335
rect 85118 262535 85174 263335
rect 87418 262535 87474 263335
rect 89626 262535 89682 263335
rect 91926 262535 91982 263335
rect 94226 262535 94282 263335
rect 96434 262535 96490 263335
rect 98734 262535 98790 263335
rect 101034 262535 101090 263335
rect 103242 262535 103298 263335
rect 105542 262535 105598 263335
rect 107842 262535 107898 263335
rect 110050 262535 110106 263335
rect 112350 262535 112406 263335
rect 114650 262535 114706 263335
rect 116950 262535 117006 263335
rect 119158 262535 119214 263335
rect 121458 262535 121514 263335
rect 123758 262535 123814 263335
rect 125966 262535 126022 263335
rect 128266 262535 128322 263335
rect 130566 262535 130622 263335
rect 132774 262535 132830 263335
rect 135074 262535 135130 263335
rect 137374 262535 137430 263335
rect 139582 262535 139638 263335
rect 141882 262535 141938 263335
rect 144182 262535 144238 263335
rect 146390 262535 146446 263335
rect 148690 262535 148746 263335
rect 150990 262535 151046 263335
rect 153290 262535 153346 263335
rect 155498 262535 155554 263335
rect 157798 262535 157854 263335
rect 160098 262535 160154 263335
rect 162306 262535 162362 263335
rect 164606 262535 164662 263335
rect 166906 262535 166962 263335
rect 169114 262535 169170 263335
rect 171414 262535 171470 263335
rect 173714 262535 173770 263335
rect 175922 262535 175978 263335
rect 178222 262535 178278 263335
rect 180522 262535 180578 263335
rect 182730 262535 182786 263335
rect 185030 262535 185086 263335
rect 187330 262535 187386 263335
rect 189630 262535 189686 263335
rect 191838 262535 191894 263335
rect 194138 262535 194194 263335
rect 196438 262535 196494 263335
rect 198646 262535 198702 263335
rect 200946 262535 201002 263335
rect 203246 262535 203302 263335
rect 205454 262535 205510 263335
rect 207754 262535 207810 263335
rect 210054 262535 210110 263335
rect 212262 262535 212318 263335
rect 214562 262535 214618 263335
rect 216862 262535 216918 263335
rect 219070 262535 219126 263335
rect 221370 262535 221426 263335
rect 223670 262535 223726 263335
rect 225970 262535 226026 263335
rect 228178 262535 228234 263335
rect 230478 262535 230534 263335
rect 232778 262535 232834 263335
rect 234986 262535 235042 263335
rect 237286 262535 237342 263335
rect 239586 262535 239642 263335
rect 241794 262535 241850 263335
rect 244094 262535 244150 263335
rect 246394 262535 246450 263335
rect 248602 262535 248658 263335
rect 250902 262535 250958 263335
rect 253202 262535 253258 263335
rect 255410 262535 255466 263335
rect 257710 262535 257766 263335
rect 260010 262535 260066 263335
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3330 0 3386 800
rect 3882 0 3938 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5446 0 5502 800
rect 5998 0 6054 800
rect 6550 0 6606 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9678 0 9734 800
rect 10230 0 10286 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12346 0 12402 800
rect 12898 0 12954 800
rect 13450 0 13506 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16118 0 16174 800
rect 16578 0 16634 800
rect 17130 0 17186 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19246 0 19302 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23478 0 23534 800
rect 24030 0 24086 800
rect 24582 0 24638 800
rect 25134 0 25190 800
rect 25594 0 25650 800
rect 26146 0 26202 800
rect 26698 0 26754 800
rect 27250 0 27306 800
rect 27802 0 27858 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29366 0 29422 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30930 0 30986 800
rect 31482 0 31538 800
rect 32034 0 32090 800
rect 32494 0 32550 800
rect 33046 0 33102 800
rect 33598 0 33654 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 37830 0 37886 800
rect 38382 0 38438 800
rect 38934 0 38990 800
rect 39486 0 39542 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 41050 0 41106 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42614 0 42670 800
rect 43166 0 43222 800
rect 43718 0 43774 800
rect 44178 0 44234 800
rect 44730 0 44786 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46386 0 46442 800
rect 46846 0 46902 800
rect 47398 0 47454 800
rect 47950 0 48006 800
rect 48502 0 48558 800
rect 48962 0 49018 800
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50618 0 50674 800
rect 51078 0 51134 800
rect 51630 0 51686 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53286 0 53342 800
rect 53746 0 53802 800
rect 54298 0 54354 800
rect 54850 0 54906 800
rect 55402 0 55458 800
rect 55862 0 55918 800
rect 56414 0 56470 800
rect 56966 0 57022 800
rect 57518 0 57574 800
rect 57978 0 58034 800
rect 58530 0 58586 800
rect 59082 0 59138 800
rect 59634 0 59690 800
rect 60186 0 60242 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62762 0 62818 800
rect 63314 0 63370 800
rect 63866 0 63922 800
rect 64418 0 64474 800
rect 64878 0 64934 800
rect 65430 0 65486 800
rect 65982 0 66038 800
rect 66534 0 66590 800
rect 67086 0 67142 800
rect 67546 0 67602 800
rect 68098 0 68154 800
rect 68650 0 68706 800
rect 69202 0 69258 800
rect 69662 0 69718 800
rect 70214 0 70270 800
rect 70766 0 70822 800
rect 71318 0 71374 800
rect 71778 0 71834 800
rect 72330 0 72386 800
rect 72882 0 72938 800
rect 73434 0 73490 800
rect 73986 0 74042 800
rect 74446 0 74502 800
rect 74998 0 75054 800
rect 75550 0 75606 800
rect 76102 0 76158 800
rect 76562 0 76618 800
rect 77114 0 77170 800
rect 77666 0 77722 800
rect 78218 0 78274 800
rect 78770 0 78826 800
rect 79230 0 79286 800
rect 79782 0 79838 800
rect 80334 0 80390 800
rect 80886 0 80942 800
rect 81346 0 81402 800
rect 81898 0 81954 800
rect 82450 0 82506 800
rect 83002 0 83058 800
rect 83462 0 83518 800
rect 84014 0 84070 800
rect 84566 0 84622 800
rect 85118 0 85174 800
rect 85670 0 85726 800
rect 86130 0 86186 800
rect 86682 0 86738 800
rect 87234 0 87290 800
rect 87786 0 87842 800
rect 88246 0 88302 800
rect 88798 0 88854 800
rect 89350 0 89406 800
rect 89902 0 89958 800
rect 90362 0 90418 800
rect 90914 0 90970 800
rect 91466 0 91522 800
rect 92018 0 92074 800
rect 92570 0 92626 800
rect 93030 0 93086 800
rect 93582 0 93638 800
rect 94134 0 94190 800
rect 94686 0 94742 800
rect 95146 0 95202 800
rect 95698 0 95754 800
rect 96250 0 96306 800
rect 96802 0 96858 800
rect 97262 0 97318 800
rect 97814 0 97870 800
rect 98366 0 98422 800
rect 98918 0 98974 800
rect 99470 0 99526 800
rect 99930 0 99986 800
rect 100482 0 100538 800
rect 101034 0 101090 800
rect 101586 0 101642 800
rect 102046 0 102102 800
rect 102598 0 102654 800
rect 103150 0 103206 800
rect 103702 0 103758 800
rect 104162 0 104218 800
rect 104714 0 104770 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106370 0 106426 800
rect 106830 0 106886 800
rect 107382 0 107438 800
rect 107934 0 107990 800
rect 108486 0 108542 800
rect 108946 0 109002 800
rect 109498 0 109554 800
rect 110050 0 110106 800
rect 110602 0 110658 800
rect 111062 0 111118 800
rect 111614 0 111670 800
rect 112166 0 112222 800
rect 112718 0 112774 800
rect 113270 0 113326 800
rect 113730 0 113786 800
rect 114282 0 114338 800
rect 114834 0 114890 800
rect 115386 0 115442 800
rect 115846 0 115902 800
rect 116398 0 116454 800
rect 116950 0 117006 800
rect 117502 0 117558 800
rect 118054 0 118110 800
rect 118514 0 118570 800
rect 119066 0 119122 800
rect 119618 0 119674 800
rect 120170 0 120226 800
rect 120630 0 120686 800
rect 121182 0 121238 800
rect 121734 0 121790 800
rect 122286 0 122342 800
rect 122746 0 122802 800
rect 123298 0 123354 800
rect 123850 0 123906 800
rect 124402 0 124458 800
rect 124954 0 125010 800
rect 125414 0 125470 800
rect 125966 0 126022 800
rect 126518 0 126574 800
rect 127070 0 127126 800
rect 127530 0 127586 800
rect 128082 0 128138 800
rect 128634 0 128690 800
rect 129186 0 129242 800
rect 129646 0 129702 800
rect 130198 0 130254 800
rect 130750 0 130806 800
rect 131302 0 131358 800
rect 131854 0 131910 800
rect 132314 0 132370 800
rect 132866 0 132922 800
rect 133418 0 133474 800
rect 133970 0 134026 800
rect 134430 0 134486 800
rect 134982 0 135038 800
rect 135534 0 135590 800
rect 136086 0 136142 800
rect 136546 0 136602 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138202 0 138258 800
rect 138754 0 138810 800
rect 139214 0 139270 800
rect 139766 0 139822 800
rect 140318 0 140374 800
rect 140870 0 140926 800
rect 141330 0 141386 800
rect 141882 0 141938 800
rect 142434 0 142490 800
rect 142986 0 143042 800
rect 143446 0 143502 800
rect 143998 0 144054 800
rect 144550 0 144606 800
rect 145102 0 145158 800
rect 145654 0 145710 800
rect 146114 0 146170 800
rect 146666 0 146722 800
rect 147218 0 147274 800
rect 147770 0 147826 800
rect 148230 0 148286 800
rect 148782 0 148838 800
rect 149334 0 149390 800
rect 149886 0 149942 800
rect 150438 0 150494 800
rect 150898 0 150954 800
rect 151450 0 151506 800
rect 152002 0 152058 800
rect 152554 0 152610 800
rect 153014 0 153070 800
rect 153566 0 153622 800
rect 154118 0 154174 800
rect 154670 0 154726 800
rect 155130 0 155186 800
rect 155682 0 155738 800
rect 156234 0 156290 800
rect 156786 0 156842 800
rect 157338 0 157394 800
rect 157798 0 157854 800
rect 158350 0 158406 800
rect 158902 0 158958 800
rect 159454 0 159510 800
rect 159914 0 159970 800
rect 160466 0 160522 800
rect 161018 0 161074 800
rect 161570 0 161626 800
rect 162030 0 162086 800
rect 162582 0 162638 800
rect 163134 0 163190 800
rect 163686 0 163742 800
rect 164238 0 164294 800
rect 164698 0 164754 800
rect 165250 0 165306 800
rect 165802 0 165858 800
rect 166354 0 166410 800
rect 166814 0 166870 800
rect 167366 0 167422 800
rect 167918 0 167974 800
rect 168470 0 168526 800
rect 168930 0 168986 800
rect 169482 0 169538 800
rect 170034 0 170090 800
rect 170586 0 170642 800
rect 171138 0 171194 800
rect 171598 0 171654 800
rect 172150 0 172206 800
rect 172702 0 172758 800
rect 173254 0 173310 800
rect 173714 0 173770 800
rect 174266 0 174322 800
rect 174818 0 174874 800
rect 175370 0 175426 800
rect 175830 0 175886 800
rect 176382 0 176438 800
rect 176934 0 176990 800
rect 177486 0 177542 800
rect 178038 0 178094 800
rect 178498 0 178554 800
rect 179050 0 179106 800
rect 179602 0 179658 800
rect 180154 0 180210 800
rect 180614 0 180670 800
rect 181166 0 181222 800
rect 181718 0 181774 800
rect 182270 0 182326 800
rect 182730 0 182786 800
rect 183282 0 183338 800
rect 183834 0 183890 800
rect 184386 0 184442 800
rect 184938 0 184994 800
rect 185398 0 185454 800
rect 185950 0 186006 800
rect 186502 0 186558 800
rect 187054 0 187110 800
rect 187514 0 187570 800
rect 188066 0 188122 800
rect 188618 0 188674 800
rect 189170 0 189226 800
rect 189722 0 189778 800
rect 190182 0 190238 800
rect 190734 0 190790 800
rect 191286 0 191342 800
rect 191838 0 191894 800
rect 192298 0 192354 800
rect 192850 0 192906 800
rect 193402 0 193458 800
rect 193954 0 194010 800
rect 194414 0 194470 800
rect 194966 0 195022 800
rect 195518 0 195574 800
rect 196070 0 196126 800
rect 196622 0 196678 800
rect 197082 0 197138 800
rect 197634 0 197690 800
rect 198186 0 198242 800
rect 198738 0 198794 800
rect 199198 0 199254 800
rect 199750 0 199806 800
rect 200302 0 200358 800
rect 200854 0 200910 800
rect 201314 0 201370 800
rect 201866 0 201922 800
rect 202418 0 202474 800
rect 202970 0 203026 800
rect 203522 0 203578 800
rect 203982 0 204038 800
rect 204534 0 204590 800
rect 205086 0 205142 800
rect 205638 0 205694 800
rect 206098 0 206154 800
rect 206650 0 206706 800
rect 207202 0 207258 800
rect 207754 0 207810 800
rect 208214 0 208270 800
rect 208766 0 208822 800
rect 209318 0 209374 800
rect 209870 0 209926 800
rect 210422 0 210478 800
rect 210882 0 210938 800
rect 211434 0 211490 800
rect 211986 0 212042 800
rect 212538 0 212594 800
rect 212998 0 213054 800
rect 213550 0 213606 800
rect 214102 0 214158 800
rect 214654 0 214710 800
rect 215114 0 215170 800
rect 215666 0 215722 800
rect 216218 0 216274 800
rect 216770 0 216826 800
rect 217322 0 217378 800
rect 217782 0 217838 800
rect 218334 0 218390 800
rect 218886 0 218942 800
rect 219438 0 219494 800
rect 219898 0 219954 800
rect 220450 0 220506 800
rect 221002 0 221058 800
rect 221554 0 221610 800
rect 222014 0 222070 800
rect 222566 0 222622 800
rect 223118 0 223174 800
rect 223670 0 223726 800
rect 224222 0 224278 800
rect 224682 0 224738 800
rect 225234 0 225290 800
rect 225786 0 225842 800
rect 226338 0 226394 800
rect 226798 0 226854 800
rect 227350 0 227406 800
rect 227902 0 227958 800
rect 228454 0 228510 800
rect 229006 0 229062 800
rect 229466 0 229522 800
rect 230018 0 230074 800
rect 230570 0 230626 800
rect 231122 0 231178 800
rect 231582 0 231638 800
rect 232134 0 232190 800
rect 232686 0 232742 800
rect 233238 0 233294 800
rect 233698 0 233754 800
rect 234250 0 234306 800
rect 234802 0 234858 800
rect 235354 0 235410 800
rect 235906 0 235962 800
rect 236366 0 236422 800
rect 236918 0 236974 800
rect 237470 0 237526 800
rect 238022 0 238078 800
rect 238482 0 238538 800
rect 239034 0 239090 800
rect 239586 0 239642 800
rect 240138 0 240194 800
rect 240598 0 240654 800
rect 241150 0 241206 800
rect 241702 0 241758 800
rect 242254 0 242310 800
rect 242806 0 242862 800
rect 243266 0 243322 800
rect 243818 0 243874 800
rect 244370 0 244426 800
rect 244922 0 244978 800
rect 245382 0 245438 800
rect 245934 0 245990 800
rect 246486 0 246542 800
rect 247038 0 247094 800
rect 247498 0 247554 800
rect 248050 0 248106 800
rect 248602 0 248658 800
rect 249154 0 249210 800
rect 249706 0 249762 800
rect 250166 0 250222 800
rect 250718 0 250774 800
rect 251270 0 251326 800
rect 251822 0 251878 800
rect 252282 0 252338 800
rect 252834 0 252890 800
rect 253386 0 253442 800
rect 253938 0 253994 800
rect 254398 0 254454 800
rect 254950 0 255006 800
rect 255502 0 255558 800
rect 256054 0 256110 800
rect 256606 0 256662 800
rect 257066 0 257122 800
rect 257618 0 257674 800
rect 258170 0 258226 800
rect 258722 0 258778 800
rect 259182 0 259238 800
rect 259734 0 259790 800
rect 260286 0 260342 800
rect 260838 0 260894 800
<< obsm2 >>
rect 204 262479 1066 262535
rect 1234 262479 3274 262535
rect 3442 262479 5574 262535
rect 5742 262479 7874 262535
rect 8042 262479 10082 262535
rect 10250 262479 12382 262535
rect 12550 262479 14682 262535
rect 14850 262479 16890 262535
rect 17058 262479 19190 262535
rect 19358 262479 21490 262535
rect 21658 262479 23698 262535
rect 23866 262479 25998 262535
rect 26166 262479 28298 262535
rect 28466 262479 30506 262535
rect 30674 262479 32806 262535
rect 32974 262479 35106 262535
rect 35274 262479 37314 262535
rect 37482 262479 39614 262535
rect 39782 262479 41914 262535
rect 42082 262479 44214 262535
rect 44382 262479 46422 262535
rect 46590 262479 48722 262535
rect 48890 262479 51022 262535
rect 51190 262479 53230 262535
rect 53398 262479 55530 262535
rect 55698 262479 57830 262535
rect 57998 262479 60038 262535
rect 60206 262479 62338 262535
rect 62506 262479 64638 262535
rect 64806 262479 66846 262535
rect 67014 262479 69146 262535
rect 69314 262479 71446 262535
rect 71614 262479 73654 262535
rect 73822 262479 75954 262535
rect 76122 262479 78254 262535
rect 78422 262479 80554 262535
rect 80722 262479 82762 262535
rect 82930 262479 85062 262535
rect 85230 262479 87362 262535
rect 87530 262479 89570 262535
rect 89738 262479 91870 262535
rect 92038 262479 94170 262535
rect 94338 262479 96378 262535
rect 96546 262479 98678 262535
rect 98846 262479 100978 262535
rect 101146 262479 103186 262535
rect 103354 262479 105486 262535
rect 105654 262479 107786 262535
rect 107954 262479 109994 262535
rect 110162 262479 112294 262535
rect 112462 262479 114594 262535
rect 114762 262479 116894 262535
rect 117062 262479 119102 262535
rect 119270 262479 121402 262535
rect 121570 262479 123702 262535
rect 123870 262479 125910 262535
rect 126078 262479 128210 262535
rect 128378 262479 130510 262535
rect 130678 262479 132718 262535
rect 132886 262479 135018 262535
rect 135186 262479 137318 262535
rect 137486 262479 139526 262535
rect 139694 262479 141826 262535
rect 141994 262479 144126 262535
rect 144294 262479 146334 262535
rect 146502 262479 148634 262535
rect 148802 262479 150934 262535
rect 151102 262479 153234 262535
rect 153402 262479 155442 262535
rect 155610 262479 157742 262535
rect 157910 262479 160042 262535
rect 160210 262479 162250 262535
rect 162418 262479 164550 262535
rect 164718 262479 166850 262535
rect 167018 262479 169058 262535
rect 169226 262479 171358 262535
rect 171526 262479 173658 262535
rect 173826 262479 175866 262535
rect 176034 262479 178166 262535
rect 178334 262479 180466 262535
rect 180634 262479 182674 262535
rect 182842 262479 184974 262535
rect 185142 262479 187274 262535
rect 187442 262479 189574 262535
rect 189742 262479 191782 262535
rect 191950 262479 194082 262535
rect 194250 262479 196382 262535
rect 196550 262479 198590 262535
rect 198758 262479 200890 262535
rect 201058 262479 203190 262535
rect 203358 262479 205398 262535
rect 205566 262479 207698 262535
rect 207866 262479 209998 262535
rect 210166 262479 212206 262535
rect 212374 262479 214506 262535
rect 214674 262479 216806 262535
rect 216974 262479 219014 262535
rect 219182 262479 221314 262535
rect 221482 262479 223614 262535
rect 223782 262479 225914 262535
rect 226082 262479 228122 262535
rect 228290 262479 230422 262535
rect 230590 262479 232722 262535
rect 232890 262479 234930 262535
rect 235098 262479 237230 262535
rect 237398 262479 239530 262535
rect 239698 262479 241738 262535
rect 241906 262479 244038 262535
rect 244206 262479 246338 262535
rect 246506 262479 248546 262535
rect 248714 262479 250846 262535
rect 251014 262479 253146 262535
rect 253314 262479 255354 262535
rect 255522 262479 257654 262535
rect 257822 262479 259954 262535
rect 260122 262479 260892 262535
rect 204 856 260892 262479
rect 314 800 606 856
rect 774 800 1158 856
rect 1326 800 1710 856
rect 1878 800 2262 856
rect 2430 800 2722 856
rect 2890 800 3274 856
rect 3442 800 3826 856
rect 3994 800 4378 856
rect 4546 800 4838 856
rect 5006 800 5390 856
rect 5558 800 5942 856
rect 6110 800 6494 856
rect 6662 800 7046 856
rect 7214 800 7506 856
rect 7674 800 8058 856
rect 8226 800 8610 856
rect 8778 800 9162 856
rect 9330 800 9622 856
rect 9790 800 10174 856
rect 10342 800 10726 856
rect 10894 800 11278 856
rect 11446 800 11738 856
rect 11906 800 12290 856
rect 12458 800 12842 856
rect 13010 800 13394 856
rect 13562 800 13946 856
rect 14114 800 14406 856
rect 14574 800 14958 856
rect 15126 800 15510 856
rect 15678 800 16062 856
rect 16230 800 16522 856
rect 16690 800 17074 856
rect 17242 800 17626 856
rect 17794 800 18178 856
rect 18346 800 18638 856
rect 18806 800 19190 856
rect 19358 800 19742 856
rect 19910 800 20294 856
rect 20462 800 20846 856
rect 21014 800 21306 856
rect 21474 800 21858 856
rect 22026 800 22410 856
rect 22578 800 22962 856
rect 23130 800 23422 856
rect 23590 800 23974 856
rect 24142 800 24526 856
rect 24694 800 25078 856
rect 25246 800 25538 856
rect 25706 800 26090 856
rect 26258 800 26642 856
rect 26810 800 27194 856
rect 27362 800 27746 856
rect 27914 800 28206 856
rect 28374 800 28758 856
rect 28926 800 29310 856
rect 29478 800 29862 856
rect 30030 800 30322 856
rect 30490 800 30874 856
rect 31042 800 31426 856
rect 31594 800 31978 856
rect 32146 800 32438 856
rect 32606 800 32990 856
rect 33158 800 33542 856
rect 33710 800 34094 856
rect 34262 800 34646 856
rect 34814 800 35106 856
rect 35274 800 35658 856
rect 35826 800 36210 856
rect 36378 800 36762 856
rect 36930 800 37222 856
rect 37390 800 37774 856
rect 37942 800 38326 856
rect 38494 800 38878 856
rect 39046 800 39430 856
rect 39598 800 39890 856
rect 40058 800 40442 856
rect 40610 800 40994 856
rect 41162 800 41546 856
rect 41714 800 42006 856
rect 42174 800 42558 856
rect 42726 800 43110 856
rect 43278 800 43662 856
rect 43830 800 44122 856
rect 44290 800 44674 856
rect 44842 800 45226 856
rect 45394 800 45778 856
rect 45946 800 46330 856
rect 46498 800 46790 856
rect 46958 800 47342 856
rect 47510 800 47894 856
rect 48062 800 48446 856
rect 48614 800 48906 856
rect 49074 800 49458 856
rect 49626 800 50010 856
rect 50178 800 50562 856
rect 50730 800 51022 856
rect 51190 800 51574 856
rect 51742 800 52126 856
rect 52294 800 52678 856
rect 52846 800 53230 856
rect 53398 800 53690 856
rect 53858 800 54242 856
rect 54410 800 54794 856
rect 54962 800 55346 856
rect 55514 800 55806 856
rect 55974 800 56358 856
rect 56526 800 56910 856
rect 57078 800 57462 856
rect 57630 800 57922 856
rect 58090 800 58474 856
rect 58642 800 59026 856
rect 59194 800 59578 856
rect 59746 800 60130 856
rect 60298 800 60590 856
rect 60758 800 61142 856
rect 61310 800 61694 856
rect 61862 800 62246 856
rect 62414 800 62706 856
rect 62874 800 63258 856
rect 63426 800 63810 856
rect 63978 800 64362 856
rect 64530 800 64822 856
rect 64990 800 65374 856
rect 65542 800 65926 856
rect 66094 800 66478 856
rect 66646 800 67030 856
rect 67198 800 67490 856
rect 67658 800 68042 856
rect 68210 800 68594 856
rect 68762 800 69146 856
rect 69314 800 69606 856
rect 69774 800 70158 856
rect 70326 800 70710 856
rect 70878 800 71262 856
rect 71430 800 71722 856
rect 71890 800 72274 856
rect 72442 800 72826 856
rect 72994 800 73378 856
rect 73546 800 73930 856
rect 74098 800 74390 856
rect 74558 800 74942 856
rect 75110 800 75494 856
rect 75662 800 76046 856
rect 76214 800 76506 856
rect 76674 800 77058 856
rect 77226 800 77610 856
rect 77778 800 78162 856
rect 78330 800 78714 856
rect 78882 800 79174 856
rect 79342 800 79726 856
rect 79894 800 80278 856
rect 80446 800 80830 856
rect 80998 800 81290 856
rect 81458 800 81842 856
rect 82010 800 82394 856
rect 82562 800 82946 856
rect 83114 800 83406 856
rect 83574 800 83958 856
rect 84126 800 84510 856
rect 84678 800 85062 856
rect 85230 800 85614 856
rect 85782 800 86074 856
rect 86242 800 86626 856
rect 86794 800 87178 856
rect 87346 800 87730 856
rect 87898 800 88190 856
rect 88358 800 88742 856
rect 88910 800 89294 856
rect 89462 800 89846 856
rect 90014 800 90306 856
rect 90474 800 90858 856
rect 91026 800 91410 856
rect 91578 800 91962 856
rect 92130 800 92514 856
rect 92682 800 92974 856
rect 93142 800 93526 856
rect 93694 800 94078 856
rect 94246 800 94630 856
rect 94798 800 95090 856
rect 95258 800 95642 856
rect 95810 800 96194 856
rect 96362 800 96746 856
rect 96914 800 97206 856
rect 97374 800 97758 856
rect 97926 800 98310 856
rect 98478 800 98862 856
rect 99030 800 99414 856
rect 99582 800 99874 856
rect 100042 800 100426 856
rect 100594 800 100978 856
rect 101146 800 101530 856
rect 101698 800 101990 856
rect 102158 800 102542 856
rect 102710 800 103094 856
rect 103262 800 103646 856
rect 103814 800 104106 856
rect 104274 800 104658 856
rect 104826 800 105210 856
rect 105378 800 105762 856
rect 105930 800 106314 856
rect 106482 800 106774 856
rect 106942 800 107326 856
rect 107494 800 107878 856
rect 108046 800 108430 856
rect 108598 800 108890 856
rect 109058 800 109442 856
rect 109610 800 109994 856
rect 110162 800 110546 856
rect 110714 800 111006 856
rect 111174 800 111558 856
rect 111726 800 112110 856
rect 112278 800 112662 856
rect 112830 800 113214 856
rect 113382 800 113674 856
rect 113842 800 114226 856
rect 114394 800 114778 856
rect 114946 800 115330 856
rect 115498 800 115790 856
rect 115958 800 116342 856
rect 116510 800 116894 856
rect 117062 800 117446 856
rect 117614 800 117998 856
rect 118166 800 118458 856
rect 118626 800 119010 856
rect 119178 800 119562 856
rect 119730 800 120114 856
rect 120282 800 120574 856
rect 120742 800 121126 856
rect 121294 800 121678 856
rect 121846 800 122230 856
rect 122398 800 122690 856
rect 122858 800 123242 856
rect 123410 800 123794 856
rect 123962 800 124346 856
rect 124514 800 124898 856
rect 125066 800 125358 856
rect 125526 800 125910 856
rect 126078 800 126462 856
rect 126630 800 127014 856
rect 127182 800 127474 856
rect 127642 800 128026 856
rect 128194 800 128578 856
rect 128746 800 129130 856
rect 129298 800 129590 856
rect 129758 800 130142 856
rect 130310 800 130694 856
rect 130862 800 131246 856
rect 131414 800 131798 856
rect 131966 800 132258 856
rect 132426 800 132810 856
rect 132978 800 133362 856
rect 133530 800 133914 856
rect 134082 800 134374 856
rect 134542 800 134926 856
rect 135094 800 135478 856
rect 135646 800 136030 856
rect 136198 800 136490 856
rect 136658 800 137042 856
rect 137210 800 137594 856
rect 137762 800 138146 856
rect 138314 800 138698 856
rect 138866 800 139158 856
rect 139326 800 139710 856
rect 139878 800 140262 856
rect 140430 800 140814 856
rect 140982 800 141274 856
rect 141442 800 141826 856
rect 141994 800 142378 856
rect 142546 800 142930 856
rect 143098 800 143390 856
rect 143558 800 143942 856
rect 144110 800 144494 856
rect 144662 800 145046 856
rect 145214 800 145598 856
rect 145766 800 146058 856
rect 146226 800 146610 856
rect 146778 800 147162 856
rect 147330 800 147714 856
rect 147882 800 148174 856
rect 148342 800 148726 856
rect 148894 800 149278 856
rect 149446 800 149830 856
rect 149998 800 150382 856
rect 150550 800 150842 856
rect 151010 800 151394 856
rect 151562 800 151946 856
rect 152114 800 152498 856
rect 152666 800 152958 856
rect 153126 800 153510 856
rect 153678 800 154062 856
rect 154230 800 154614 856
rect 154782 800 155074 856
rect 155242 800 155626 856
rect 155794 800 156178 856
rect 156346 800 156730 856
rect 156898 800 157282 856
rect 157450 800 157742 856
rect 157910 800 158294 856
rect 158462 800 158846 856
rect 159014 800 159398 856
rect 159566 800 159858 856
rect 160026 800 160410 856
rect 160578 800 160962 856
rect 161130 800 161514 856
rect 161682 800 161974 856
rect 162142 800 162526 856
rect 162694 800 163078 856
rect 163246 800 163630 856
rect 163798 800 164182 856
rect 164350 800 164642 856
rect 164810 800 165194 856
rect 165362 800 165746 856
rect 165914 800 166298 856
rect 166466 800 166758 856
rect 166926 800 167310 856
rect 167478 800 167862 856
rect 168030 800 168414 856
rect 168582 800 168874 856
rect 169042 800 169426 856
rect 169594 800 169978 856
rect 170146 800 170530 856
rect 170698 800 171082 856
rect 171250 800 171542 856
rect 171710 800 172094 856
rect 172262 800 172646 856
rect 172814 800 173198 856
rect 173366 800 173658 856
rect 173826 800 174210 856
rect 174378 800 174762 856
rect 174930 800 175314 856
rect 175482 800 175774 856
rect 175942 800 176326 856
rect 176494 800 176878 856
rect 177046 800 177430 856
rect 177598 800 177982 856
rect 178150 800 178442 856
rect 178610 800 178994 856
rect 179162 800 179546 856
rect 179714 800 180098 856
rect 180266 800 180558 856
rect 180726 800 181110 856
rect 181278 800 181662 856
rect 181830 800 182214 856
rect 182382 800 182674 856
rect 182842 800 183226 856
rect 183394 800 183778 856
rect 183946 800 184330 856
rect 184498 800 184882 856
rect 185050 800 185342 856
rect 185510 800 185894 856
rect 186062 800 186446 856
rect 186614 800 186998 856
rect 187166 800 187458 856
rect 187626 800 188010 856
rect 188178 800 188562 856
rect 188730 800 189114 856
rect 189282 800 189666 856
rect 189834 800 190126 856
rect 190294 800 190678 856
rect 190846 800 191230 856
rect 191398 800 191782 856
rect 191950 800 192242 856
rect 192410 800 192794 856
rect 192962 800 193346 856
rect 193514 800 193898 856
rect 194066 800 194358 856
rect 194526 800 194910 856
rect 195078 800 195462 856
rect 195630 800 196014 856
rect 196182 800 196566 856
rect 196734 800 197026 856
rect 197194 800 197578 856
rect 197746 800 198130 856
rect 198298 800 198682 856
rect 198850 800 199142 856
rect 199310 800 199694 856
rect 199862 800 200246 856
rect 200414 800 200798 856
rect 200966 800 201258 856
rect 201426 800 201810 856
rect 201978 800 202362 856
rect 202530 800 202914 856
rect 203082 800 203466 856
rect 203634 800 203926 856
rect 204094 800 204478 856
rect 204646 800 205030 856
rect 205198 800 205582 856
rect 205750 800 206042 856
rect 206210 800 206594 856
rect 206762 800 207146 856
rect 207314 800 207698 856
rect 207866 800 208158 856
rect 208326 800 208710 856
rect 208878 800 209262 856
rect 209430 800 209814 856
rect 209982 800 210366 856
rect 210534 800 210826 856
rect 210994 800 211378 856
rect 211546 800 211930 856
rect 212098 800 212482 856
rect 212650 800 212942 856
rect 213110 800 213494 856
rect 213662 800 214046 856
rect 214214 800 214598 856
rect 214766 800 215058 856
rect 215226 800 215610 856
rect 215778 800 216162 856
rect 216330 800 216714 856
rect 216882 800 217266 856
rect 217434 800 217726 856
rect 217894 800 218278 856
rect 218446 800 218830 856
rect 218998 800 219382 856
rect 219550 800 219842 856
rect 220010 800 220394 856
rect 220562 800 220946 856
rect 221114 800 221498 856
rect 221666 800 221958 856
rect 222126 800 222510 856
rect 222678 800 223062 856
rect 223230 800 223614 856
rect 223782 800 224166 856
rect 224334 800 224626 856
rect 224794 800 225178 856
rect 225346 800 225730 856
rect 225898 800 226282 856
rect 226450 800 226742 856
rect 226910 800 227294 856
rect 227462 800 227846 856
rect 228014 800 228398 856
rect 228566 800 228950 856
rect 229118 800 229410 856
rect 229578 800 229962 856
rect 230130 800 230514 856
rect 230682 800 231066 856
rect 231234 800 231526 856
rect 231694 800 232078 856
rect 232246 800 232630 856
rect 232798 800 233182 856
rect 233350 800 233642 856
rect 233810 800 234194 856
rect 234362 800 234746 856
rect 234914 800 235298 856
rect 235466 800 235850 856
rect 236018 800 236310 856
rect 236478 800 236862 856
rect 237030 800 237414 856
rect 237582 800 237966 856
rect 238134 800 238426 856
rect 238594 800 238978 856
rect 239146 800 239530 856
rect 239698 800 240082 856
rect 240250 800 240542 856
rect 240710 800 241094 856
rect 241262 800 241646 856
rect 241814 800 242198 856
rect 242366 800 242750 856
rect 242918 800 243210 856
rect 243378 800 243762 856
rect 243930 800 244314 856
rect 244482 800 244866 856
rect 245034 800 245326 856
rect 245494 800 245878 856
rect 246046 800 246430 856
rect 246598 800 246982 856
rect 247150 800 247442 856
rect 247610 800 247994 856
rect 248162 800 248546 856
rect 248714 800 249098 856
rect 249266 800 249650 856
rect 249818 800 250110 856
rect 250278 800 250662 856
rect 250830 800 251214 856
rect 251382 800 251766 856
rect 251934 800 252226 856
rect 252394 800 252778 856
rect 252946 800 253330 856
rect 253498 800 253882 856
rect 254050 800 254342 856
rect 254510 800 254894 856
rect 255062 800 255446 856
rect 255614 800 255998 856
rect 256166 800 256550 856
rect 256718 800 257010 856
rect 257178 800 257562 856
rect 257730 800 258114 856
rect 258282 800 258666 856
rect 258834 800 259126 856
rect 259294 800 259678 856
rect 259846 800 260230 856
rect 260398 800 260782 856
<< obsm3 >>
rect 2865 1939 253907 261153
<< metal4 >>
rect 4208 2128 4528 261168
rect 4868 2176 5188 261120
rect 5528 2176 5848 261120
rect 6188 2176 6508 261120
rect 19568 2128 19888 261168
rect 20228 2176 20548 261120
rect 20888 2176 21208 261120
rect 21548 2176 21868 261120
rect 34928 2128 35248 261168
rect 35588 2176 35908 261120
rect 36248 2176 36568 261120
rect 36908 2176 37228 261120
rect 50288 2128 50608 261168
rect 50948 2176 51268 261120
rect 51608 2176 51928 261120
rect 52268 2176 52588 261120
rect 65648 2128 65968 261168
rect 66308 2176 66628 261120
rect 66968 2176 67288 261120
rect 67628 2176 67948 261120
rect 81008 2128 81328 261168
rect 81668 2176 81988 261120
rect 82328 2176 82648 261120
rect 82988 2176 83308 261120
rect 96368 2128 96688 261168
rect 97028 2176 97348 261120
rect 97688 2176 98008 261120
rect 98348 2176 98668 261120
rect 111728 2128 112048 261168
rect 112388 2176 112708 261120
rect 113048 2176 113368 261120
rect 113708 2176 114028 261120
rect 127088 2128 127408 261168
rect 127748 2176 128068 261120
rect 128408 2176 128728 261120
rect 129068 2176 129388 261120
rect 142448 2128 142768 261168
rect 143108 2176 143428 261120
rect 143768 2176 144088 261120
rect 144428 2176 144748 261120
rect 157808 2128 158128 261168
rect 158468 2176 158788 261120
rect 159128 2176 159448 261120
rect 159788 2176 160108 261120
rect 173168 2128 173488 261168
rect 173828 2176 174148 261120
rect 174488 2176 174808 261120
rect 175148 2176 175468 261120
rect 188528 2128 188848 261168
rect 189188 2176 189508 261120
rect 189848 2176 190168 261120
rect 190508 2176 190828 261120
rect 203888 2128 204208 261168
rect 204548 2176 204868 261120
rect 205208 2176 205528 261120
rect 205868 2176 206188 261120
rect 219248 2128 219568 261168
rect 219908 2176 220228 261120
rect 220568 2176 220888 261120
rect 221228 2176 221548 261120
rect 234608 2128 234928 261168
rect 235268 2176 235588 261120
rect 235928 2176 236248 261120
rect 236588 2176 236908 261120
rect 249968 2128 250288 261168
rect 250628 2176 250948 261120
rect 251288 2176 251608 261120
rect 251948 2176 252268 261120
<< obsm4 >>
rect 50107 57835 50208 239597
rect 50688 57835 50868 239597
rect 51348 57835 51528 239597
rect 52008 57835 52188 239597
rect 52668 57835 65568 239597
rect 66048 57835 66228 239597
rect 66708 57835 66888 239597
rect 67368 57835 67548 239597
rect 68028 57835 80928 239597
rect 81408 57835 81588 239597
rect 82068 57835 82248 239597
rect 82728 57835 82908 239597
rect 83388 57835 96288 239597
rect 96768 57835 96948 239597
rect 97428 57835 97608 239597
rect 98088 57835 98268 239597
rect 98748 57835 111648 239597
rect 112128 57835 112308 239597
rect 112788 57835 112968 239597
rect 113448 57835 113628 239597
rect 114108 57835 127008 239597
rect 127488 57835 127668 239597
rect 128148 57835 128328 239597
rect 128808 57835 128988 239597
rect 129468 57835 142368 239597
rect 142848 57835 143028 239597
rect 143508 57835 143688 239597
rect 144168 57835 144348 239597
rect 144828 57835 157728 239597
rect 158208 57835 158388 239597
rect 158868 57835 159048 239597
rect 159528 57835 159708 239597
rect 160188 57835 173088 239597
rect 173568 57835 173748 239597
rect 174228 57835 174408 239597
rect 174888 57835 175068 239597
rect 175548 57835 188448 239597
rect 188928 57835 189108 239597
rect 189588 57835 189768 239597
rect 190248 57835 190428 239597
rect 190908 57835 203808 239597
rect 204288 57835 204468 239597
rect 204948 57835 205128 239597
rect 205608 57835 205788 239597
rect 206268 57835 219168 239597
rect 219648 57835 219828 239597
rect 220308 57835 220488 239597
rect 220968 57835 221148 239597
rect 221628 57835 234528 239597
rect 235008 57835 235093 239597
<< labels >>
rlabel metal2 s 1122 262535 1178 263335 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 69202 262535 69258 263335 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 76010 262535 76066 263335 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 82818 262535 82874 263335 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 89626 262535 89682 263335 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 96434 262535 96490 263335 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 103242 262535 103298 263335 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 110050 262535 110106 263335 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 116950 262535 117006 263335 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 123758 262535 123814 263335 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 130566 262535 130622 263335 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7930 262535 7986 263335 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 137374 262535 137430 263335 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 144182 262535 144238 263335 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 150990 262535 151046 263335 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 157798 262535 157854 263335 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 164606 262535 164662 263335 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 171414 262535 171470 263335 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 178222 262535 178278 263335 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 185030 262535 185086 263335 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 191838 262535 191894 263335 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 198646 262535 198702 263335 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14738 262535 14794 263335 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 205454 262535 205510 263335 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 212262 262535 212318 263335 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 219070 262535 219126 263335 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 225970 262535 226026 263335 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 232778 262535 232834 263335 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 239586 262535 239642 263335 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 246394 262535 246450 263335 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 253202 262535 253258 263335 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 21546 262535 21602 263335 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 28354 262535 28410 263335 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 35162 262535 35218 263335 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 41970 262535 42026 263335 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 48778 262535 48834 263335 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 55586 262535 55642 263335 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 62394 262535 62450 263335 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3330 262535 3386 263335 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 71502 262535 71558 263335 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 78310 262535 78366 263335 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 85118 262535 85174 263335 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 91926 262535 91982 263335 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 98734 262535 98790 263335 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 105542 262535 105598 263335 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 112350 262535 112406 263335 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 119158 262535 119214 263335 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 125966 262535 126022 263335 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 132774 262535 132830 263335 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 10138 262535 10194 263335 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 139582 262535 139638 263335 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 146390 262535 146446 263335 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 153290 262535 153346 263335 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 160098 262535 160154 263335 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 166906 262535 166962 263335 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 173714 262535 173770 263335 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 180522 262535 180578 263335 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 187330 262535 187386 263335 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 194138 262535 194194 263335 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 200946 262535 201002 263335 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 16946 262535 17002 263335 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 207754 262535 207810 263335 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 214562 262535 214618 263335 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 221370 262535 221426 263335 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 228178 262535 228234 263335 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 234986 262535 235042 263335 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 241794 262535 241850 263335 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 248602 262535 248658 263335 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 255410 262535 255466 263335 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 23754 262535 23810 263335 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 30562 262535 30618 263335 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 37370 262535 37426 263335 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 44270 262535 44326 263335 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 51078 262535 51134 263335 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 57886 262535 57942 263335 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 64694 262535 64750 263335 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5630 262535 5686 263335 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 73710 262535 73766 263335 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 80610 262535 80666 263335 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 87418 262535 87474 263335 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 94226 262535 94282 263335 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 101034 262535 101090 263335 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 107842 262535 107898 263335 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 114650 262535 114706 263335 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 121458 262535 121514 263335 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 128266 262535 128322 263335 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 135074 262535 135130 263335 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 12438 262535 12494 263335 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 141882 262535 141938 263335 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 148690 262535 148746 263335 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 155498 262535 155554 263335 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 162306 262535 162362 263335 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 169114 262535 169170 263335 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 175922 262535 175978 263335 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 182730 262535 182786 263335 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 189630 262535 189686 263335 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 196438 262535 196494 263335 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 203246 262535 203302 263335 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 19246 262535 19302 263335 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 210054 262535 210110 263335 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 216862 262535 216918 263335 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 223670 262535 223726 263335 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 230478 262535 230534 263335 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 237286 262535 237342 263335 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 244094 262535 244150 263335 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 250902 262535 250958 263335 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 257710 262535 257766 263335 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 26054 262535 26110 263335 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 32862 262535 32918 263335 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 39670 262535 39726 263335 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 46478 262535 46534 263335 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 53286 262535 53342 263335 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 60094 262535 60150 263335 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 66902 262535 66958 263335 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 260010 262535 260066 263335 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 260286 0 260342 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 260838 0 260894 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 218886 0 218942 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 222014 0 222070 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 223670 0 223726 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 225234 0 225290 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 239586 0 239642 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 241150 0 241206 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 242806 0 242862 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 244370 0 244426 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 245934 0 245990 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 247498 0 247554 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 249154 0 249210 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 250718 0 250774 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 252282 0 252338 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 255502 0 255558 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 257066 0 257122 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 258722 0 258778 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 187054 0 187110 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 191838 0 191894 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 193402 0 193458 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 198186 0 198242 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 201314 0 201370 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 202970 0 203026 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 207754 0 207810 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 214102 0 214158 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 216218 0 216274 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 217782 0 217838 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 219438 0 219494 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 221002 0 221058 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 222566 0 222622 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 225786 0 225842 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 227350 0 227406 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 229006 0 229062 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 230570 0 230626 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 232134 0 232190 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 233698 0 233754 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 235354 0 235410 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 236918 0 236974 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 238482 0 238538 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 240138 0 240194 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 241702 0 241758 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 243266 0 243322 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 244922 0 244978 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 246486 0 246542 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 248050 0 248106 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 249706 0 249762 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 251270 0 251326 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 252834 0 252890 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 254398 0 254454 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 256054 0 256110 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 257618 0 257674 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 259182 0 259238 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 131854 0 131910 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 141330 0 141386 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 155682 0 155738 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 163686 0 163742 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 165250 0 165306 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 168470 0 168526 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 176382 0 176438 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 179602 0 179658 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 181166 0 181222 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 182730 0 182786 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 184386 0 184442 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 187514 0 187570 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 189170 0 189226 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 190734 0 190790 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 193954 0 194010 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 195518 0 195574 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 198738 0 198794 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 200302 0 200358 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 201866 0 201922 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 203522 0 203578 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 205086 0 205142 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 206650 0 206706 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 208214 0 208270 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 209870 0 209926 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 211434 0 211490 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 212998 0 213054 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 214654 0 214710 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 216770 0 216826 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 224682 0 224738 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 227902 0 227958 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 229466 0 229522 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 232686 0 232742 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 234250 0 234306 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 235906 0 235962 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 237470 0 237526 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 240598 0 240654 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 242254 0 242310 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 243818 0 243874 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 251822 0 251878 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 254950 0 255006 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 256606 0 256662 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 258170 0 258226 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 259734 0 259790 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 186502 0 186558 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 202418 0 202474 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 203982 0 204038 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 208766 0 208822 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 213550 0 213606 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 249968 2128 250288 261168 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 261168 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 261168 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 261168 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 261168 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 261168 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 261168 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 261168 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 261168 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 234608 2128 234928 261168 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 261168 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 261168 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 261168 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 261168 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 261168 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 261168 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 261168 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 250628 2176 250948 261120 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 261120 6 vccd2
port 626 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 261120 6 vccd2
port 627 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 261120 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 261120 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 261120 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 261120 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 261120 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 261120 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 235268 2176 235588 261120 6 vssd2
port 634 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 261120 6 vssd2
port 635 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 261120 6 vssd2
port 636 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 261120 6 vssd2
port 637 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 261120 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 261120 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 261120 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 261120 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 251288 2176 251608 261120 6 vdda1
port 642 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 261120 6 vdda1
port 643 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 261120 6 vdda1
port 644 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 261120 6 vdda1
port 645 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 261120 6 vdda1
port 646 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 261120 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 261120 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 261120 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 261120 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 235928 2176 236248 261120 6 vssa1
port 651 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 261120 6 vssa1
port 652 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 261120 6 vssa1
port 653 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 261120 6 vssa1
port 654 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 261120 6 vssa1
port 655 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 261120 6 vssa1
port 656 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 261120 6 vssa1
port 657 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 261120 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 251948 2176 252268 261120 6 vdda2
port 659 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 261120 6 vdda2
port 660 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 261120 6 vdda2
port 661 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 261120 6 vdda2
port 662 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 261120 6 vdda2
port 663 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 261120 6 vdda2
port 664 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 261120 6 vdda2
port 665 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 261120 6 vdda2
port 666 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 261120 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 236588 2176 236908 261120 6 vssa2
port 668 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 261120 6 vssa2
port 669 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 261120 6 vssa2
port 670 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 261120 6 vssa2
port 671 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 261120 6 vssa2
port 672 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 261120 6 vssa2
port 673 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 261120 6 vssa2
port 674 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 261120 6 vssa2
port 675 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 261191 263335
string LEFview TRUE
string GDS_FILE /project/openlane/axi_dma/runs/axi_dma/results/magic/axi_dma.gds
string GDS_END 95171696
string GDS_START 1124848
<< end >>

